* Example HSPICE testbench file (test.sp)
* transistor model
.INCLUDE "/cae/apps/data/asap7PDK-2022/asap7PDK_r1p7/models/hspice/7nm_TT_160803.pm"

* Design Under Test (DUT)
.INCLUDE "Neuron.sp" * Enable this line for schematic netlist

*.INCLUDE "INV.pex.netlist" * Enable this line for layout netlist
* Simulation Parameters
.TEMP 25.0
.options artist=2 ingold=2 parhier=local psf=2 hier_delim=0 accurate=1 NUMDGT=8 measdgt=5 GMINDC=1e-18 DELMAX=1n method=gear INGOLD=2 POST=1

.subckt INV_V2 a vdd vss y
mn0 y a vss vss nmos_rvt w=54e-9 l=20e-9 nfin=1
mp1 y a vdd vdd pmos_rvt w=81e-9 l=20e-9 nfin=1
.ends INV_V2

xi24 z0<0> vdd vss inv_out INV_V2
xi23 z0<0> vdd vss inv_out INV_V2
xi22 z0<0> vdd vss inv_out2 INV_V2
xi21 z0<0> vdd vss inv_out INV_V2
xi28 z0<1> vdd vss inv_out INV_V2
xi27 z0<1> vdd vss inv_out INV_V2
xi26 z0<1> vdd vss inv_out2 INV_V2
xi25 z0<1> vdd vss inv_out INV_V2

* Instantiate (DUT)
xd1  VDD VSS  W01<1> X1<0> W00<1> X0<0> X1<1> W01<0> X0<1> W00<0> 
+ W20<0> W20<1> W20<2> 
+ Z0<1> Z0<0> 
+ Neuron
vdd0 vdd vss 0.9v
vss0 vss 0 0v

V_X0<1> X0<1> 0 PWL(0.000000n 0.0  0.100000n 0.0  0.125000n 0.0  0.225000n 0.0  0.250000n 0.0  0.350000n 0.0  0.375000n 0.0  0.475000n 0.0  0.500000n 0.0  0.600000n 0.0  0.625000n 0.0  0.725000n 0.0  0.750000n 0.0  0.850000n 0.0  0.875000n 0.0  0.975000n 0.0  1.000000n 0.0  1.100000n 0.0  1.125000n 0.0  1.225000n 0.0  1.250000n 0.0  1.350000n 0.0  1.375000n 0.0  1.475000n 0.0  1.500000n 0.0  1.600000n 0.0  1.625000n 0.0  1.725000n 0.0  1.750000n 0.0  1.850000n 0.0  1.875000n 0.0  1.975000n 0.0  2.000000n 0.0  2.100000n 0.0  2.125000n 0.0  2.225000n 0.0  2.250000n 0.0  2.350000n 0.0  2.375000n 0.0  2.475000n 0.0  2.500000n 0.0  2.600000n 0.0  2.625000n 0.0  2.725000n 0.0  2.750000n 0.0  2.850000n 0.0  2.875000n 0.0  2.975000n 0.0  3.000000n 0.0  3.100000n 0.0  3.125000n 0.0  3.225000n 0.0  3.250000n 0.0  3.350000n 0.0  3.375000n 0.0  3.475000n 0.0  3.500000n 0.0  3.600000n 0.0  3.625000n 0.0  3.725000n 0.0  3.750000n 0.0  3.850000n 0.0  3.875000n 0.0  3.975000n 0.0  4.000000n 0.0  4.100000n 0.0  4.125000n 0.0  4.225000n 0.0  4.250000n 0.0  4.350000n 0.0  4.375000n 0.0  4.475000n 0.0  4.500000n 0.0  4.600000n 0.0  4.625000n 0.0  4.725000n 0.0  4.750000n 0.0  4.850000n 0.0  4.875000n 0.0  4.975000n 0.0  5.000000n 0.0  5.100000n 0.0  5.125000n 0.0  5.225000n 0.0  5.250000n 0.0  5.350000n 0.0  5.375000n 0.0  5.475000n 0.0  5.500000n 0.0  5.600000n 0.0  5.625000n 0.0  5.725000n 0.0  5.750000n 0.0  5.850000n 0.0  5.875000n 0.0  5.975000n 0.0  6.000000n 0.0  6.100000n 0.0  6.125000n 0.0  6.225000n 0.0  6.250000n 0.0  6.350000n 0.0  6.375000n 0.0  6.475000n 0.0  6.500000n 0.0  6.600000n 0.0  6.625000n 0.0  6.725000n 0.0  6.750000n 0.0  6.850000n 0.0  6.875000n 0.0  6.975000n 0.0  7.000000n 0.0  7.100000n 0.0  7.125000n 0.0  7.225000n 0.0  7.250000n 0.0  7.350000n 0.0  7.375000n 0.0  7.475000n 0.0  7.500000n 0.0  7.600000n 0.0  7.625000n 0.0  7.725000n 0.0  7.750000n 0.0  7.850000n 0.0  7.875000n 0.0  7.975000n 0.0  8.000000n 0.0  8.100000n 0.0  8.125000n 0.0  8.225000n 0.0  8.250000n 0.0  8.350000n 0.0  8.375000n 0.0  8.475000n 0.0  8.500000n 0.0  8.600000n 0.0  8.625000n 0.0  8.725000n 0.0  8.750000n 0.0  8.850000n 0.0  8.875000n 0.0  8.975000n 0.0  9.000000n 0.0  9.100000n 0.0  9.125000n 0.0  9.225000n 0.0  9.250000n 0.0  9.350000n 0.0  9.375000n 0.0  9.475000n 0.0  9.500000n 0.0  9.600000n 0.0  9.625000n 0.0  9.725000n 0.0  9.750000n 0.0  9.850000n 0.0  9.875000n 0.0  9.975000n 0.0  10.000000n 0.0  10.100000n 0.0  10.125000n 0.0  10.225000n 0.0  10.250000n 0.0  10.350000n 0.0  10.375000n 0.0  10.475000n 0.0  10.500000n 0.0  10.600000n 0.0  10.625000n 0.0  10.725000n 0.0  10.750000n 0.0  10.850000n 0.0  10.875000n 0.0  10.975000n 0.0  11.000000n 0.0  11.100000n 0.0  11.125000n 0.0  11.225000n 0.0  11.250000n 0.0  11.350000n 0.0  11.375000n 0.0  11.475000n 0.0  11.500000n 0.0  11.600000n 0.0  11.625000n 0.0  11.725000n 0.0  11.750000n 0.0  11.850000n 0.0  11.875000n 0.0  11.975000n 0.0  12.000000n 0.0  12.100000n 0.0  12.125000n 0.0  12.225000n 0.0  12.250000n 0.0  12.350000n 0.0  12.375000n 0.0  12.475000n 0.0  12.500000n 0.0  12.600000n 0.0  12.625000n 0.0  12.725000n 0.0  12.750000n 0.0  12.850000n 0.0  12.875000n 0.0  12.975000n 0.0  13.000000n 0.0  13.100000n 0.0  13.125000n 0.0  13.225000n 0.0  13.250000n 0.0  13.350000n 0.0  13.375000n 0.0  13.475000n 0.0  13.500000n 0.0  13.600000n 0.0  13.625000n 0.0  13.725000n 0.0  13.750000n 0.0  13.850000n 0.0  13.875000n 0.0  13.975000n 0.0  14.000000n 0.0  14.100000n 0.0  14.125000n 0.0  14.225000n 0.0  14.250000n 0.0  14.350000n 0.0  14.375000n 0.0  14.475000n 0.0  14.500000n 0.0  14.600000n 0.0  14.625000n 0.0  14.725000n 0.0  14.750000n 0.0  14.850000n 0.0  14.875000n 0.0  14.975000n 0.0  15.000000n 0.0  15.100000n 0.0  15.125000n 0.0  15.225000n 0.0  15.250000n 0.0  15.350000n 0.0  15.375000n 0.0  15.475000n 0.0  15.500000n 0.0  15.600000n 0.0  15.625000n 0.0  15.725000n 0.0  15.750000n 0.0  15.850000n 0.0  15.875000n 0.0  15.975000n 0.0  16.000000n 0.0  16.100000n 0.0  16.125000n 0.0  16.225000n 0.0  16.250000n 0.0  16.350000n 0.0  16.375000n 0.0  16.475000n 0.0  16.500000n 0.0  16.600000n 0.0  16.625000n 0.0  16.725000n 0.0  16.750000n 0.0  16.850000n 0.0  16.875000n 0.0  16.975000n 0.0  17.000000n 0.0  17.100000n 0.0  17.125000n 0.0  17.225000n 0.0  17.250000n 0.0  17.350000n 0.0  17.375000n 0.0  17.475000n 0.0  17.500000n 0.0  17.600000n 0.0  17.625000n 0.0  17.725000n 0.0  17.750000n 0.0  17.850000n 0.0  17.875000n 0.0  17.975000n 0.0  18.000000n 0.0  18.100000n 0.0  18.125000n 0.0  18.225000n 0.0  18.250000n 0.0  18.350000n 0.0  18.375000n 0.0  18.475000n 0.0  18.500000n 0.0  18.600000n 0.0  18.625000n 0.0  18.725000n 0.0  18.750000n 0.0  18.850000n 0.0  18.875000n 0.0  18.975000n 0.0  19.000000n 0.0  19.100000n 0.0  19.125000n 0.0  19.225000n 0.0  19.250000n 0.0  19.350000n 0.0  19.375000n 0.0  19.475000n 0.0  19.500000n 0.0  19.600000n 0.0  19.625000n 0.0  19.725000n 0.0  19.750000n 0.0  19.850000n 0.0  19.875000n 0.0  19.975000n 0.0  20.000000n 0.0  20.100000n 0.0  20.125000n 0.0  20.225000n 0.0  20.250000n 0.9  20.350000n 0.9  20.375000n 0.9  20.475000n 0.9  20.500000n 0.9  20.600000n 0.9  20.625000n 0.9  20.725000n 0.9  20.750000n 0.9  20.850000n 0.9  20.875000n 0.9  20.975000n 0.9  21.000000n 0.9  21.100000n 0.9  21.125000n 0.9  21.225000n 0.9  21.250000n 0.9  21.350000n 0.9  21.375000n 0.9  21.475000n 0.9  21.500000n 0.9  21.600000n 0.9  21.625000n 0.9  21.725000n 0.9  21.750000n 0.9  21.850000n 0.9  21.875000n 0.9  21.975000n 0.9  22.000000n 0.9  22.100000n 0.9  22.125000n 0.9  22.225000n 0.9  22.250000n 0.9  22.350000n 0.9  22.375000n 0.9  22.475000n 0.9  22.500000n 0.9  22.600000n 0.9  22.625000n 0.9  22.725000n 0.9  22.750000n 0.9  22.850000n 0.9  22.875000n 0.9  22.975000n 0.9  23.000000n 0.9  23.100000n 0.9  23.125000n 0.9  23.225000n 0.9  23.250000n 0.9  23.350000n 0.9  23.375000n 0.9  23.475000n 0.9  23.500000n 0.9  23.600000n 0.9  23.625000n 0.9  23.725000n 0.9  23.750000n 0.9  23.850000n 0.9  23.875000n 0.9  23.975000n 0.9  24.000000n 0.9  24.100000n 0.9  24.125000n 0.9  24.225000n 0.9  24.250000n 0.9  24.350000n 0.9  24.375000n 0.9  24.475000n 0.9  24.500000n 0.9  24.600000n 0.9  24.625000n 0.9  24.725000n 0.9  24.750000n 0.9  24.850000n 0.9  24.875000n 0.9  24.975000n 0.9  25.000000n 0.9  25.100000n 0.9  25.125000n 0.9  25.225000n 0.9  25.250000n 0.9  25.350000n 0.9  25.375000n 0.9  25.475000n 0.9  25.500000n 0.9  25.600000n 0.9  25.625000n 0.9  25.725000n 0.9  25.750000n 0.9  25.850000n 0.9  25.875000n 0.9  25.975000n 0.9  26.000000n 0.9  26.100000n 0.9  26.125000n 0.9  26.225000n 0.9  26.250000n 0.9  26.350000n 0.9  26.375000n 0.9  26.475000n 0.9  26.500000n 0.9  26.600000n 0.9  26.625000n 0.9  26.725000n 0.9  26.750000n 0.9  26.850000n 0.9  26.875000n 0.9  26.975000n 0.9  27.000000n 0.9  27.100000n 0.9  27.125000n 0.9  27.225000n 0.9  27.250000n 0.9  27.350000n 0.9  27.375000n 0.9  27.475000n 0.9  27.500000n 0.9  27.600000n 0.9  27.625000n 0.9  27.725000n 0.9  27.750000n 0.9  27.850000n 0.9  27.875000n 0.9  27.975000n 0.9  28.000000n 0.9  28.100000n 0.9  28.125000n 0.9  28.225000n 0.9  28.250000n 0.9  28.350000n 0.9  28.375000n 0.9  28.475000n 0.9  28.500000n 0.9  28.600000n 0.9  28.625000n 0.9  28.725000n 0.9  28.750000n 0.9  28.850000n 0.9  28.875000n 0.9  28.975000n 0.9  29.000000n 0.9  29.100000n 0.9  29.125000n 0.9  29.225000n 0.9  29.250000n 0.9  29.350000n 0.9  29.375000n 0.9  29.475000n 0.9  29.500000n 0.9  29.600000n 0.9  29.625000n 0.9  29.725000n 0.9  29.750000n 0.9  29.850000n 0.9  29.875000n 0.9  29.975000n 0.9  30.000000n 0.9  30.100000n 0.9  30.125000n 0.9  30.225000n 0.9  30.250000n 0.9 )
V_X0<0> X0<0> 0 PWL(0.000000n 0.0  0.100000n 0.0  0.125000n 0.0  0.225000n 0.0  0.250000n 0.0  0.350000n 0.0  0.375000n 0.0  0.475000n 0.0  0.500000n 0.0  0.600000n 0.0  0.625000n 0.0  0.725000n 0.0  0.750000n 0.0  0.850000n 0.0  0.875000n 0.0  0.975000n 0.0  1.000000n 0.0  1.100000n 0.0  1.125000n 0.0  1.225000n 0.0  1.250000n 0.0  1.350000n 0.0  1.375000n 0.0  1.475000n 0.0  1.500000n 0.0  1.600000n 0.0  1.625000n 0.0  1.725000n 0.0  1.750000n 0.0  1.850000n 0.0  1.875000n 0.0  1.975000n 0.0  2.000000n 0.0  2.100000n 0.0  2.125000n 0.0  2.225000n 0.0  2.250000n 0.0  2.350000n 0.0  2.375000n 0.0  2.475000n 0.0  2.500000n 0.0  2.600000n 0.0  2.625000n 0.0  2.725000n 0.0  2.750000n 0.0  2.850000n 0.0  2.875000n 0.0  2.975000n 0.0  3.000000n 0.0  3.100000n 0.0  3.125000n 0.0  3.225000n 0.0  3.250000n 0.0  3.350000n 0.0  3.375000n 0.0  3.475000n 0.0  3.500000n 0.0  3.600000n 0.0  3.625000n 0.0  3.725000n 0.0  3.750000n 0.0  3.850000n 0.0  3.875000n 0.0  3.975000n 0.0  4.000000n 0.0  4.100000n 0.0  4.125000n 0.0  4.225000n 0.0  4.250000n 0.0  4.350000n 0.0  4.375000n 0.0  4.475000n 0.0  4.500000n 0.0  4.600000n 0.0  4.625000n 0.0  4.725000n 0.0  4.750000n 0.0  4.850000n 0.0  4.875000n 0.0  4.975000n 0.0  5.000000n 0.0  5.100000n 0.0  5.125000n 0.0  5.225000n 0.0  5.250000n 0.0  5.350000n 0.0  5.375000n 0.0  5.475000n 0.0  5.500000n 0.0  5.600000n 0.0  5.625000n 0.0  5.725000n 0.0  5.750000n 0.0  5.850000n 0.0  5.875000n 0.0  5.975000n 0.0  6.000000n 0.0  6.100000n 0.0  6.125000n 0.0  6.225000n 0.0  6.250000n 0.0  6.350000n 0.0  6.375000n 0.0  6.475000n 0.0  6.500000n 0.0  6.600000n 0.0  6.625000n 0.0  6.725000n 0.0  6.750000n 0.0  6.850000n 0.0  6.875000n 0.0  6.975000n 0.0  7.000000n 0.0  7.100000n 0.0  7.125000n 0.0  7.225000n 0.0  7.250000n 0.0  7.350000n 0.0  7.375000n 0.0  7.475000n 0.0  7.500000n 0.0  7.600000n 0.0  7.625000n 0.0  7.725000n 0.0  7.750000n 0.0  7.850000n 0.0  7.875000n 0.0  7.975000n 0.0  8.000000n 0.0  8.100000n 0.0  8.125000n 0.0  8.225000n 0.0  8.250000n 0.0  8.350000n 0.0  8.375000n 0.0  8.475000n 0.0  8.500000n 0.0  8.600000n 0.0  8.625000n 0.0  8.725000n 0.0  8.750000n 0.0  8.850000n 0.0  8.875000n 0.0  8.975000n 0.0  9.000000n 0.0  9.100000n 0.0  9.125000n 0.0  9.225000n 0.0  9.250000n 0.0  9.350000n 0.0  9.375000n 0.0  9.475000n 0.0  9.500000n 0.0  9.600000n 0.0  9.625000n 0.0  9.725000n 0.0  9.750000n 0.0  9.850000n 0.0  9.875000n 0.0  9.975000n 0.0  10.000000n 0.0  10.100000n 0.0  10.125000n 0.9  10.225000n 0.9  10.250000n 0.9  10.350000n 0.9  10.375000n 0.9  10.475000n 0.9  10.500000n 0.9  10.600000n 0.9  10.625000n 0.9  10.725000n 0.9  10.750000n 0.9  10.850000n 0.9  10.875000n 0.9  10.975000n 0.9  11.000000n 0.9  11.100000n 0.9  11.125000n 0.9  11.225000n 0.9  11.250000n 0.9  11.350000n 0.9  11.375000n 0.9  11.475000n 0.9  11.500000n 0.9  11.600000n 0.9  11.625000n 0.9  11.725000n 0.9  11.750000n 0.9  11.850000n 0.9  11.875000n 0.9  11.975000n 0.9  12.000000n 0.9  12.100000n 0.9  12.125000n 0.9  12.225000n 0.9  12.250000n 0.9  12.350000n 0.9  12.375000n 0.9  12.475000n 0.9  12.500000n 0.9  12.600000n 0.9  12.625000n 0.9  12.725000n 0.9  12.750000n 0.9  12.850000n 0.9  12.875000n 0.9  12.975000n 0.9  13.000000n 0.9  13.100000n 0.9  13.125000n 0.9  13.225000n 0.9  13.250000n 0.9  13.350000n 0.9  13.375000n 0.9  13.475000n 0.9  13.500000n 0.9  13.600000n 0.9  13.625000n 0.9  13.725000n 0.9  13.750000n 0.9  13.850000n 0.9  13.875000n 0.9  13.975000n 0.9  14.000000n 0.9  14.100000n 0.9  14.125000n 0.9  14.225000n 0.9  14.250000n 0.9  14.350000n 0.9  14.375000n 0.9  14.475000n 0.9  14.500000n 0.9  14.600000n 0.9  14.625000n 0.9  14.725000n 0.9  14.750000n 0.9  14.850000n 0.9  14.875000n 0.9  14.975000n 0.9  15.000000n 0.9  15.100000n 0.9  15.125000n 0.9  15.225000n 0.9  15.250000n 0.9  15.350000n 0.9  15.375000n 0.9  15.475000n 0.9  15.500000n 0.9  15.600000n 0.9  15.625000n 0.9  15.725000n 0.9  15.750000n 0.9  15.850000n 0.9  15.875000n 0.9  15.975000n 0.9  16.000000n 0.9  16.100000n 0.9  16.125000n 0.9  16.225000n 0.9  16.250000n 0.9  16.350000n 0.9  16.375000n 0.9  16.475000n 0.9  16.500000n 0.9  16.600000n 0.9  16.625000n 0.9  16.725000n 0.9  16.750000n 0.9  16.850000n 0.9  16.875000n 0.9  16.975000n 0.9  17.000000n 0.9  17.100000n 0.9  17.125000n 0.9  17.225000n 0.9  17.250000n 0.9  17.350000n 0.9  17.375000n 0.9  17.475000n 0.9  17.500000n 0.9  17.600000n 0.9  17.625000n 0.9  17.725000n 0.9  17.750000n 0.9  17.850000n 0.9  17.875000n 0.9  17.975000n 0.9  18.000000n 0.9  18.100000n 0.9  18.125000n 0.9  18.225000n 0.9  18.250000n 0.9  18.350000n 0.9  18.375000n 0.9  18.475000n 0.9  18.500000n 0.9  18.600000n 0.9  18.625000n 0.9  18.725000n 0.9  18.750000n 0.9  18.850000n 0.9  18.875000n 0.9  18.975000n 0.9  19.000000n 0.9  19.100000n 0.9  19.125000n 0.9  19.225000n 0.9  19.250000n 0.9  19.350000n 0.9  19.375000n 0.9  19.475000n 0.9  19.500000n 0.9  19.600000n 0.9  19.625000n 0.9  19.725000n 0.9  19.750000n 0.9  19.850000n 0.9  19.875000n 0.9  19.975000n 0.9  20.000000n 0.9  20.100000n 0.9  20.125000n 0.9  20.225000n 0.9  20.250000n 0.9  20.350000n 0.9  20.375000n 0.9  20.475000n 0.9  20.500000n 0.9  20.600000n 0.9  20.625000n 0.9  20.725000n 0.9  20.750000n 0.9  20.850000n 0.9  20.875000n 0.9  20.975000n 0.9  21.000000n 0.9  21.100000n 0.9  21.125000n 0.9  21.225000n 0.9  21.250000n 0.9  21.350000n 0.9  21.375000n 0.9  21.475000n 0.9  21.500000n 0.9  21.600000n 0.9  21.625000n 0.9  21.725000n 0.9  21.750000n 0.9  21.850000n 0.9  21.875000n 0.9  21.975000n 0.9  22.000000n 0.9  22.100000n 0.9  22.125000n 0.9  22.225000n 0.9  22.250000n 0.9  22.350000n 0.9  22.375000n 0.9  22.475000n 0.9  22.500000n 0.9  22.600000n 0.9  22.625000n 0.9  22.725000n 0.9  22.750000n 0.9  22.850000n 0.9  22.875000n 0.9  22.975000n 0.9  23.000000n 0.9  23.100000n 0.9  23.125000n 0.9  23.225000n 0.9  23.250000n 0.9  23.350000n 0.9  23.375000n 0.9  23.475000n 0.9  23.500000n 0.9  23.600000n 0.9  23.625000n 0.9  23.725000n 0.9  23.750000n 0.9  23.850000n 0.9  23.875000n 0.9  23.975000n 0.9  24.000000n 0.9  24.100000n 0.9  24.125000n 0.9  24.225000n 0.9  24.250000n 0.9  24.350000n 0.9  24.375000n 0.9  24.475000n 0.9  24.500000n 0.9  24.600000n 0.9  24.625000n 0.9  24.725000n 0.9  24.750000n 0.9  24.850000n 0.9  24.875000n 0.9  24.975000n 0.9  25.000000n 0.9  25.100000n 0.9  25.125000n 0.9  25.225000n 0.9  25.250000n 0.9  25.350000n 0.9  25.375000n 0.9  25.475000n 0.9  25.500000n 0.9  25.600000n 0.9  25.625000n 0.9  25.725000n 0.9  25.750000n 0.9  25.850000n 0.9  25.875000n 0.9  25.975000n 0.9  26.000000n 0.9  26.100000n 0.9  26.125000n 0.9  26.225000n 0.9  26.250000n 0.9  26.350000n 0.9  26.375000n 0.9  26.475000n 0.9  26.500000n 0.9  26.600000n 0.9  26.625000n 0.9  26.725000n 0.9  26.750000n 0.9  26.850000n 0.9  26.875000n 0.9  26.975000n 0.9  27.000000n 0.9  27.100000n 0.9  27.125000n 0.9  27.225000n 0.9  27.250000n 0.9  27.350000n 0.9  27.375000n 0.9  27.475000n 0.9  27.500000n 0.9  27.600000n 0.9  27.625000n 0.9  27.725000n 0.9  27.750000n 0.9  27.850000n 0.9  27.875000n 0.9  27.975000n 0.9  28.000000n 0.9  28.100000n 0.9  28.125000n 0.9  28.225000n 0.9  28.250000n 0.9  28.350000n 0.9  28.375000n 0.9  28.475000n 0.9  28.500000n 0.9  28.600000n 0.9  28.625000n 0.9  28.725000n 0.9  28.750000n 0.9  28.850000n 0.9  28.875000n 0.9  28.975000n 0.9  29.000000n 0.9  29.100000n 0.9  29.125000n 0.9  29.225000n 0.9  29.250000n 0.9  29.350000n 0.9  29.375000n 0.9  29.475000n 0.9  29.500000n 0.9  29.600000n 0.9  29.625000n 0.9  29.725000n 0.9  29.750000n 0.9  29.850000n 0.9  29.875000n 0.9  29.975000n 0.9  30.000000n 0.9  30.100000n 0.9  30.125000n 0.9  30.225000n 0.9  30.250000n 0.9 )
V_X1<1> X1<1> 0 PWL(0.000000n 0.0  0.100000n 0.0  0.125000n 0.0  0.225000n 0.0  0.250000n 0.0  0.350000n 0.0  0.375000n 0.0  0.475000n 0.0  0.500000n 0.0  0.600000n 0.0  0.625000n 0.0  0.725000n 0.0  0.750000n 0.0  0.850000n 0.0  0.875000n 0.0  0.975000n 0.0  1.000000n 0.0  1.100000n 0.0  1.125000n 0.0  1.225000n 0.0  1.250000n 0.0  1.350000n 0.0  1.375000n 0.0  1.475000n 0.0  1.500000n 0.0  1.600000n 0.0  1.625000n 0.0  1.725000n 0.0  1.750000n 0.0  1.850000n 0.0  1.875000n 0.0  1.975000n 0.0  2.000000n 0.0  2.100000n 0.0  2.125000n 0.0  2.225000n 0.0  2.250000n 0.0  2.350000n 0.0  2.375000n 0.0  2.475000n 0.0  2.500000n 0.0  2.600000n 0.0  2.625000n 0.0  2.725000n 0.0  2.750000n 0.0  2.850000n 0.0  2.875000n 0.0  2.975000n 0.0  3.000000n 0.0  3.100000n 0.0  3.125000n 0.0  3.225000n 0.0  3.250000n 0.0  3.350000n 0.0  3.375000n 0.0  3.475000n 0.0  3.500000n 0.0  3.600000n 0.0  3.625000n 0.0  3.725000n 0.0  3.750000n 0.0  3.850000n 0.0  3.875000n 0.0  3.975000n 0.0  4.000000n 0.0  4.100000n 0.0  4.125000n 0.0  4.225000n 0.0  4.250000n 0.0  4.350000n 0.0  4.375000n 0.0  4.475000n 0.0  4.500000n 0.0  4.600000n 0.0  4.625000n 0.0  4.725000n 0.0  4.750000n 0.0  4.850000n 0.0  4.875000n 0.0  4.975000n 0.0  5.000000n 0.0  5.100000n 0.0  5.125000n 0.0  5.225000n 0.0  5.250000n 0.0  5.350000n 0.0  5.375000n 0.0  5.475000n 0.0  5.500000n 0.0  5.600000n 0.0  5.625000n 0.0  5.725000n 0.0  5.750000n 0.0  5.850000n 0.0  5.875000n 0.0  5.975000n 0.0  6.000000n 0.0  6.100000n 0.0  6.125000n 0.0  6.225000n 0.0  6.250000n 0.0  6.350000n 0.0  6.375000n 0.0  6.475000n 0.0  6.500000n 0.0  6.600000n 0.0  6.625000n 0.0  6.725000n 0.0  6.750000n 0.9  6.850000n 0.9  6.875000n 0.9  6.975000n 0.9  7.000000n 0.9  7.100000n 0.9  7.125000n 0.9  7.225000n 0.9  7.250000n 0.9  7.350000n 0.9  7.375000n 0.9  7.475000n 0.9  7.500000n 0.9  7.600000n 0.9  7.625000n 0.9  7.725000n 0.9  7.750000n 0.9  7.850000n 0.9  7.875000n 0.9  7.975000n 0.9  8.000000n 0.9  8.100000n 0.9  8.125000n 0.9  8.225000n 0.9  8.250000n 0.9  8.350000n 0.9  8.375000n 0.9  8.475000n 0.9  8.500000n 0.9  8.600000n 0.9  8.625000n 0.9  8.725000n 0.9  8.750000n 0.9  8.850000n 0.9  8.875000n 0.9  8.975000n 0.9  9.000000n 0.9  9.100000n 0.9  9.125000n 0.9  9.225000n 0.9  9.250000n 0.9  9.350000n 0.9  9.375000n 0.9  9.475000n 0.9  9.500000n 0.9  9.600000n 0.9  9.625000n 0.9  9.725000n 0.9  9.750000n 0.9  9.850000n 0.9  9.875000n 0.9  9.975000n 0.9  10.000000n 0.9  10.100000n 0.9  10.125000n 0.9  10.225000n 0.9  10.250000n 0.9  10.350000n 0.9  10.375000n 0.9  10.475000n 0.9  10.500000n 0.9  10.600000n 0.9  10.625000n 0.9  10.725000n 0.9  10.750000n 0.9  10.850000n 0.9  10.875000n 0.9  10.975000n 0.9  11.000000n 0.9  11.100000n 0.9  11.125000n 0.9  11.225000n 0.9  11.250000n 0.9  11.350000n 0.9  11.375000n 0.9  11.475000n 0.9  11.500000n 0.9  11.600000n 0.9  11.625000n 0.9  11.725000n 0.9  11.750000n 0.9  11.850000n 0.9  11.875000n 0.9  11.975000n 0.9  12.000000n 0.9  12.100000n 0.9  12.125000n 0.9  12.225000n 0.9  12.250000n 0.9  12.350000n 0.9  12.375000n 0.9  12.475000n 0.9  12.500000n 0.9  12.600000n 0.9  12.625000n 0.9  12.725000n 0.9  12.750000n 0.9  12.850000n 0.9  12.875000n 0.9  12.975000n 0.9  13.000000n 0.9  13.100000n 0.9  13.125000n 0.9  13.225000n 0.9  13.250000n 0.9  13.350000n 0.9  13.375000n 0.9  13.475000n 0.9  13.500000n 0.0  13.600000n 0.0  13.625000n 0.0  13.725000n 0.0  13.750000n 0.0  13.850000n 0.0  13.875000n 0.0  13.975000n 0.0  14.000000n 0.0  14.100000n 0.0  14.125000n 0.0  14.225000n 0.0  14.250000n 0.0  14.350000n 0.0  14.375000n 0.0  14.475000n 0.0  14.500000n 0.0  14.600000n 0.0  14.625000n 0.0  14.725000n 0.0  14.750000n 0.0  14.850000n 0.0  14.875000n 0.0  14.975000n 0.0  15.000000n 0.0  15.100000n 0.0  15.125000n 0.0  15.225000n 0.0  15.250000n 0.0  15.350000n 0.0  15.375000n 0.0  15.475000n 0.0  15.500000n 0.0  15.600000n 0.0  15.625000n 0.0  15.725000n 0.0  15.750000n 0.0  15.850000n 0.0  15.875000n 0.0  15.975000n 0.0  16.000000n 0.0  16.100000n 0.0  16.125000n 0.0  16.225000n 0.0  16.250000n 0.0  16.350000n 0.0  16.375000n 0.0  16.475000n 0.0  16.500000n 0.0  16.600000n 0.0  16.625000n 0.0  16.725000n 0.0  16.750000n 0.0  16.850000n 0.0  16.875000n 0.0  16.975000n 0.0  17.000000n 0.0  17.100000n 0.0  17.125000n 0.0  17.225000n 0.0  17.250000n 0.0  17.350000n 0.0  17.375000n 0.0  17.475000n 0.0  17.500000n 0.0  17.600000n 0.0  17.625000n 0.0  17.725000n 0.0  17.750000n 0.0  17.850000n 0.0  17.875000n 0.0  17.975000n 0.0  18.000000n 0.0  18.100000n 0.0  18.125000n 0.0  18.225000n 0.0  18.250000n 0.0  18.350000n 0.0  18.375000n 0.0  18.475000n 0.0  18.500000n 0.0  18.600000n 0.0  18.625000n 0.0  18.725000n 0.0  18.750000n 0.0  18.850000n 0.0  18.875000n 0.0  18.975000n 0.0  19.000000n 0.0  19.100000n 0.0  19.125000n 0.0  19.225000n 0.0  19.250000n 0.0  19.350000n 0.0  19.375000n 0.0  19.475000n 0.0  19.500000n 0.0  19.600000n 0.0  19.625000n 0.0  19.725000n 0.0  19.750000n 0.0  19.850000n 0.0  19.875000n 0.0  19.975000n 0.0  20.000000n 0.0  20.100000n 0.0  20.125000n 0.0  20.225000n 0.0  20.250000n 0.0  20.350000n 0.0  20.375000n 0.0  20.475000n 0.0  20.500000n 0.0  20.600000n 0.0  20.625000n 0.0  20.725000n 0.0  20.750000n 0.0  20.850000n 0.0  20.875000n 0.0  20.975000n 0.0  21.000000n 0.0  21.100000n 0.0  21.125000n 0.0  21.225000n 0.0  21.250000n 0.0  21.350000n 0.0  21.375000n 0.0  21.475000n 0.0  21.500000n 0.0  21.600000n 0.0  21.625000n 0.0  21.725000n 0.0  21.750000n 0.0  21.850000n 0.0  21.875000n 0.0  21.975000n 0.0  22.000000n 0.0  22.100000n 0.0  22.125000n 0.0  22.225000n 0.0  22.250000n 0.0  22.350000n 0.0  22.375000n 0.0  22.475000n 0.0  22.500000n 0.0  22.600000n 0.0  22.625000n 0.0  22.725000n 0.0  22.750000n 0.0  22.850000n 0.0  22.875000n 0.0  22.975000n 0.0  23.000000n 0.0  23.100000n 0.0  23.125000n 0.0  23.225000n 0.0  23.250000n 0.0  23.350000n 0.0  23.375000n 0.0  23.475000n 0.0  23.500000n 0.0  23.600000n 0.0  23.625000n 0.0  23.725000n 0.0  23.750000n 0.0  23.850000n 0.0  23.875000n 0.0  23.975000n 0.0  24.000000n 0.0  24.100000n 0.0  24.125000n 0.0  24.225000n 0.0  24.250000n 0.0  24.350000n 0.0  24.375000n 0.0  24.475000n 0.0  24.500000n 0.0  24.600000n 0.0  24.625000n 0.0  24.725000n 0.0  24.750000n 0.0  24.850000n 0.0  24.875000n 0.0  24.975000n 0.0  25.000000n 0.0  25.100000n 0.0  25.125000n 0.0  25.225000n 0.0  25.250000n 0.0  25.350000n 0.0  25.375000n 0.0  25.475000n 0.0  25.500000n 0.0  25.600000n 0.0  25.625000n 0.0  25.725000n 0.0  25.750000n 0.0  25.850000n 0.0  25.875000n 0.0  25.975000n 0.0  26.000000n 0.0  26.100000n 0.0  26.125000n 0.0  26.225000n 0.0  26.250000n 0.0  26.350000n 0.0  26.375000n 0.0  26.475000n 0.0  26.500000n 0.0  26.600000n 0.0  26.625000n 0.0  26.725000n 0.0  26.750000n 0.0  26.850000n 0.0  26.875000n 0.0  26.975000n 0.0  27.000000n 0.9  27.100000n 0.9  27.125000n 0.9  27.225000n 0.9  27.250000n 0.9  27.350000n 0.9  27.375000n 0.9  27.475000n 0.9  27.500000n 0.9  27.600000n 0.9  27.625000n 0.9  27.725000n 0.9  27.750000n 0.9  27.850000n 0.9  27.875000n 0.9  27.975000n 0.9  28.000000n 0.9  28.100000n 0.9  28.125000n 0.9  28.225000n 0.9  28.250000n 0.9  28.350000n 0.9  28.375000n 0.9  28.475000n 0.9  28.500000n 0.9  28.600000n 0.9  28.625000n 0.9  28.725000n 0.9  28.750000n 0.9  28.850000n 0.9  28.875000n 0.9  28.975000n 0.9  29.000000n 0.9  29.100000n 0.9  29.125000n 0.9  29.225000n 0.9  29.250000n 0.9  29.350000n 0.9  29.375000n 0.9  29.475000n 0.9  29.500000n 0.9  29.600000n 0.9  29.625000n 0.9  29.725000n 0.9  29.750000n 0.9  29.850000n 0.9  29.875000n 0.9  29.975000n 0.9  30.000000n 0.9  30.100000n 0.9  30.125000n 0.9  30.225000n 0.9  30.250000n 0.9 )
V_X1<0> X1<0> 0 PWL(0.000000n 0.0  0.100000n 0.0  0.125000n 0.0  0.225000n 0.0  0.250000n 0.0  0.350000n 0.0  0.375000n 0.0  0.475000n 0.0  0.500000n 0.0  0.600000n 0.0  0.625000n 0.0  0.725000n 0.0  0.750000n 0.0  0.850000n 0.0  0.875000n 0.0  0.975000n 0.0  1.000000n 0.0  1.100000n 0.0  1.125000n 0.0  1.225000n 0.0  1.250000n 0.0  1.350000n 0.0  1.375000n 0.0  1.475000n 0.0  1.500000n 0.0  1.600000n 0.0  1.625000n 0.0  1.725000n 0.0  1.750000n 0.0  1.850000n 0.0  1.875000n 0.0  1.975000n 0.0  2.000000n 0.0  2.100000n 0.0  2.125000n 0.0  2.225000n 0.0  2.250000n 0.0  2.350000n 0.0  2.375000n 0.0  2.475000n 0.0  2.500000n 0.0  2.600000n 0.0  2.625000n 0.0  2.725000n 0.0  2.750000n 0.0  2.850000n 0.0  2.875000n 0.0  2.975000n 0.0  3.000000n 0.0  3.100000n 0.0  3.125000n 0.0  3.225000n 0.0  3.250000n 0.0  3.350000n 0.0  3.375000n 0.9  3.475000n 0.9  3.500000n 0.9  3.600000n 0.9  3.625000n 0.9  3.725000n 0.9  3.750000n 0.9  3.850000n 0.9  3.875000n 0.9  3.975000n 0.9  4.000000n 0.9  4.100000n 0.9  4.125000n 0.9  4.225000n 0.9  4.250000n 0.9  4.350000n 0.9  4.375000n 0.9  4.475000n 0.9  4.500000n 0.9  4.600000n 0.9  4.625000n 0.9  4.725000n 0.9  4.750000n 0.9  4.850000n 0.9  4.875000n 0.9  4.975000n 0.9  5.000000n 0.9  5.100000n 0.9  5.125000n 0.9  5.225000n 0.9  5.250000n 0.9  5.350000n 0.9  5.375000n 0.9  5.475000n 0.9  5.500000n 0.9  5.600000n 0.9  5.625000n 0.9  5.725000n 0.9  5.750000n 0.9  5.850000n 0.9  5.875000n 0.9  5.975000n 0.9  6.000000n 0.9  6.100000n 0.9  6.125000n 0.9  6.225000n 0.9  6.250000n 0.9  6.350000n 0.9  6.375000n 0.9  6.475000n 0.9  6.500000n 0.9  6.600000n 0.9  6.625000n 0.9  6.725000n 0.9  6.750000n 0.9  6.850000n 0.9  6.875000n 0.9  6.975000n 0.9  7.000000n 0.9  7.100000n 0.9  7.125000n 0.9  7.225000n 0.9  7.250000n 0.9  7.350000n 0.9  7.375000n 0.9  7.475000n 0.9  7.500000n 0.9  7.600000n 0.9  7.625000n 0.9  7.725000n 0.9  7.750000n 0.9  7.850000n 0.9  7.875000n 0.9  7.975000n 0.9  8.000000n 0.9  8.100000n 0.9  8.125000n 0.9  8.225000n 0.9  8.250000n 0.9  8.350000n 0.9  8.375000n 0.9  8.475000n 0.9  8.500000n 0.9  8.600000n 0.9  8.625000n 0.9  8.725000n 0.9  8.750000n 0.9  8.850000n 0.9  8.875000n 0.9  8.975000n 0.9  9.000000n 0.9  9.100000n 0.9  9.125000n 0.9  9.225000n 0.9  9.250000n 0.9  9.350000n 0.9  9.375000n 0.9  9.475000n 0.9  9.500000n 0.9  9.600000n 0.9  9.625000n 0.9  9.725000n 0.9  9.750000n 0.9  9.850000n 0.9  9.875000n 0.9  9.975000n 0.9  10.000000n 0.9  10.100000n 0.9  10.125000n 0.9  10.225000n 0.9  10.250000n 0.9  10.350000n 0.9  10.375000n 0.9  10.475000n 0.9  10.500000n 0.9  10.600000n 0.9  10.625000n 0.9  10.725000n 0.9  10.750000n 0.9  10.850000n 0.9  10.875000n 0.9  10.975000n 0.9  11.000000n 0.9  11.100000n 0.9  11.125000n 0.9  11.225000n 0.9  11.250000n 0.9  11.350000n 0.9  11.375000n 0.9  11.475000n 0.9  11.500000n 0.9  11.600000n 0.9  11.625000n 0.9  11.725000n 0.9  11.750000n 0.9  11.850000n 0.9  11.875000n 0.9  11.975000n 0.9  12.000000n 0.9  12.100000n 0.9  12.125000n 0.9  12.225000n 0.9  12.250000n 0.9  12.350000n 0.9  12.375000n 0.9  12.475000n 0.9  12.500000n 0.9  12.600000n 0.9  12.625000n 0.9  12.725000n 0.9  12.750000n 0.9  12.850000n 0.9  12.875000n 0.9  12.975000n 0.9  13.000000n 0.9  13.100000n 0.9  13.125000n 0.9  13.225000n 0.9  13.250000n 0.9  13.350000n 0.9  13.375000n 0.9  13.475000n 0.9  13.500000n 0.9  13.600000n 0.9  13.625000n 0.9  13.725000n 0.9  13.750000n 0.9  13.850000n 0.9  13.875000n 0.9  13.975000n 0.9  14.000000n 0.9  14.100000n 0.9  14.125000n 0.9  14.225000n 0.9  14.250000n 0.9  14.350000n 0.9  14.375000n 0.9  14.475000n 0.9  14.500000n 0.9  14.600000n 0.9  14.625000n 0.9  14.725000n 0.9  14.750000n 0.9  14.850000n 0.9  14.875000n 0.9  14.975000n 0.9  15.000000n 0.9  15.100000n 0.9  15.125000n 0.9  15.225000n 0.9  15.250000n 0.9  15.350000n 0.9  15.375000n 0.9  15.475000n 0.9  15.500000n 0.9  15.600000n 0.9  15.625000n 0.9  15.725000n 0.9  15.750000n 0.9  15.850000n 0.9  15.875000n 0.9  15.975000n 0.9  16.000000n 0.9  16.100000n 0.9  16.125000n 0.9  16.225000n 0.9  16.250000n 0.9  16.350000n 0.9  16.375000n 0.9  16.475000n 0.9  16.500000n 0.9  16.600000n 0.9  16.625000n 0.9  16.725000n 0.9  16.750000n 0.9  16.850000n 0.9  16.875000n 0.0  16.975000n 0.0  17.000000n 0.0  17.100000n 0.0  17.125000n 0.0  17.225000n 0.0  17.250000n 0.0  17.350000n 0.0  17.375000n 0.0  17.475000n 0.0  17.500000n 0.0  17.600000n 0.0  17.625000n 0.0  17.725000n 0.0  17.750000n 0.0  17.850000n 0.0  17.875000n 0.0  17.975000n 0.0  18.000000n 0.0  18.100000n 0.0  18.125000n 0.0  18.225000n 0.0  18.250000n 0.0  18.350000n 0.0  18.375000n 0.0  18.475000n 0.0  18.500000n 0.0  18.600000n 0.0  18.625000n 0.0  18.725000n 0.0  18.750000n 0.0  18.850000n 0.0  18.875000n 0.0  18.975000n 0.0  19.000000n 0.0  19.100000n 0.0  19.125000n 0.0  19.225000n 0.0  19.250000n 0.0  19.350000n 0.0  19.375000n 0.0  19.475000n 0.0  19.500000n 0.0  19.600000n 0.0  19.625000n 0.0  19.725000n 0.0  19.750000n 0.0  19.850000n 0.0  19.875000n 0.0  19.975000n 0.0  20.000000n 0.0  20.100000n 0.0  20.125000n 0.0  20.225000n 0.0  20.250000n 0.0  20.350000n 0.0  20.375000n 0.0  20.475000n 0.0  20.500000n 0.0  20.600000n 0.0  20.625000n 0.0  20.725000n 0.0  20.750000n 0.0  20.850000n 0.0  20.875000n 0.0  20.975000n 0.0  21.000000n 0.0  21.100000n 0.0  21.125000n 0.0  21.225000n 0.0  21.250000n 0.0  21.350000n 0.0  21.375000n 0.0  21.475000n 0.0  21.500000n 0.0  21.600000n 0.0  21.625000n 0.0  21.725000n 0.0  21.750000n 0.0  21.850000n 0.0  21.875000n 0.0  21.975000n 0.0  22.000000n 0.0  22.100000n 0.0  22.125000n 0.0  22.225000n 0.0  22.250000n 0.0  22.350000n 0.0  22.375000n 0.0  22.475000n 0.0  22.500000n 0.0  22.600000n 0.0  22.625000n 0.0  22.725000n 0.0  22.750000n 0.0  22.850000n 0.0  22.875000n 0.0  22.975000n 0.0  23.000000n 0.0  23.100000n 0.0  23.125000n 0.0  23.225000n 0.0  23.250000n 0.0  23.350000n 0.0  23.375000n 0.0  23.475000n 0.0  23.500000n 0.0  23.600000n 0.0  23.625000n 0.9  23.725000n 0.9  23.750000n 0.9  23.850000n 0.9  23.875000n 0.9  23.975000n 0.9  24.000000n 0.9  24.100000n 0.9  24.125000n 0.9  24.225000n 0.9  24.250000n 0.9  24.350000n 0.9  24.375000n 0.9  24.475000n 0.9  24.500000n 0.9  24.600000n 0.9  24.625000n 0.9  24.725000n 0.9  24.750000n 0.9  24.850000n 0.9  24.875000n 0.9  24.975000n 0.9  25.000000n 0.9  25.100000n 0.9  25.125000n 0.9  25.225000n 0.9  25.250000n 0.9  25.350000n 0.9  25.375000n 0.9  25.475000n 0.9  25.500000n 0.9  25.600000n 0.9  25.625000n 0.9  25.725000n 0.9  25.750000n 0.9  25.850000n 0.9  25.875000n 0.9  25.975000n 0.9  26.000000n 0.9  26.100000n 0.9  26.125000n 0.9  26.225000n 0.9  26.250000n 0.9  26.350000n 0.9  26.375000n 0.9  26.475000n 0.9  26.500000n 0.9  26.600000n 0.9  26.625000n 0.9  26.725000n 0.9  26.750000n 0.9  26.850000n 0.9  26.875000n 0.9  26.975000n 0.9  27.000000n 0.9  27.100000n 0.9  27.125000n 0.9  27.225000n 0.9  27.250000n 0.9  27.350000n 0.9  27.375000n 0.9  27.475000n 0.9  27.500000n 0.9  27.600000n 0.9  27.625000n 0.9  27.725000n 0.9  27.750000n 0.9  27.850000n 0.9  27.875000n 0.9  27.975000n 0.9  28.000000n 0.9  28.100000n 0.9  28.125000n 0.9  28.225000n 0.9  28.250000n 0.9  28.350000n 0.9  28.375000n 0.9  28.475000n 0.9  28.500000n 0.9  28.600000n 0.9  28.625000n 0.9  28.725000n 0.9  28.750000n 0.9  28.850000n 0.9  28.875000n 0.9  28.975000n 0.9  29.000000n 0.9  29.100000n 0.9  29.125000n 0.9  29.225000n 0.9  29.250000n 0.9  29.350000n 0.9  29.375000n 0.9  29.475000n 0.9  29.500000n 0.9  29.600000n 0.9  29.625000n 0.9  29.725000n 0.9  29.750000n 0.9  29.850000n 0.9  29.875000n 0.9  29.975000n 0.9  30.000000n 0.9  30.100000n 0.9  30.125000n 0.9  30.225000n 0.9  30.250000n 0.9 )
V_W00<1> W00<1> 0 PWL(0.000000n 0.0  0.100000n 0.0  0.125000n 0.0  0.225000n 0.0  0.250000n 0.0  0.350000n 0.0  0.375000n 0.0  0.475000n 0.0  0.500000n 0.0  0.600000n 0.0  0.625000n 0.0  0.725000n 0.0  0.750000n 0.0  0.850000n 0.0  0.875000n 0.0  0.975000n 0.0  1.000000n 0.0  1.100000n 0.0  1.125000n 0.0  1.225000n 0.0  1.250000n 0.0  1.350000n 0.0  1.375000n 0.0  1.475000n 0.0  1.500000n 0.0  1.600000n 0.0  1.625000n 0.0  1.725000n 0.0  1.750000n 0.0  1.850000n 0.0  1.875000n 0.0  1.975000n 0.0  2.000000n 0.0  2.100000n 0.0  2.125000n 0.0  2.225000n 0.0  2.250000n 0.9  2.350000n 0.9  2.375000n 0.9  2.475000n 0.9  2.500000n 0.9  2.600000n 0.9  2.625000n 0.9  2.725000n 0.9  2.750000n 0.9  2.850000n 0.9  2.875000n 0.9  2.975000n 0.9  3.000000n 0.9  3.100000n 0.9  3.125000n 0.9  3.225000n 0.9  3.250000n 0.9  3.350000n 0.9  3.375000n 0.9  3.475000n 0.9  3.500000n 0.9  3.600000n 0.9  3.625000n 0.9  3.725000n 0.9  3.750000n 0.9  3.850000n 0.9  3.875000n 0.9  3.975000n 0.9  4.000000n 0.9  4.100000n 0.9  4.125000n 0.9  4.225000n 0.9  4.250000n 0.9  4.350000n 0.9  4.375000n 0.9  4.475000n 0.9  4.500000n 0.0  4.600000n 0.0  4.625000n 0.0  4.725000n 0.0  4.750000n 0.0  4.850000n 0.0  4.875000n 0.0  4.975000n 0.0  5.000000n 0.0  5.100000n 0.0  5.125000n 0.0  5.225000n 0.0  5.250000n 0.0  5.350000n 0.0  5.375000n 0.0  5.475000n 0.0  5.500000n 0.0  5.600000n 0.0  5.625000n 0.0  5.725000n 0.0  5.750000n 0.0  5.850000n 0.0  5.875000n 0.0  5.975000n 0.0  6.000000n 0.0  6.100000n 0.0  6.125000n 0.0  6.225000n 0.0  6.250000n 0.0  6.350000n 0.0  6.375000n 0.0  6.475000n 0.0  6.500000n 0.0  6.600000n 0.0  6.625000n 0.0  6.725000n 0.0  6.750000n 0.0  6.850000n 0.0  6.875000n 0.0  6.975000n 0.0  7.000000n 0.0  7.100000n 0.0  7.125000n 0.0  7.225000n 0.0  7.250000n 0.0  7.350000n 0.0  7.375000n 0.0  7.475000n 0.0  7.500000n 0.0  7.600000n 0.0  7.625000n 0.0  7.725000n 0.0  7.750000n 0.0  7.850000n 0.0  7.875000n 0.0  7.975000n 0.0  8.000000n 0.0  8.100000n 0.0  8.125000n 0.0  8.225000n 0.0  8.250000n 0.0  8.350000n 0.0  8.375000n 0.0  8.475000n 0.0  8.500000n 0.0  8.600000n 0.0  8.625000n 0.0  8.725000n 0.0  8.750000n 0.0  8.850000n 0.0  8.875000n 0.0  8.975000n 0.0  9.000000n 0.9  9.100000n 0.9  9.125000n 0.9  9.225000n 0.9  9.250000n 0.9  9.350000n 0.9  9.375000n 0.9  9.475000n 0.9  9.500000n 0.9  9.600000n 0.9  9.625000n 0.9  9.725000n 0.9  9.750000n 0.9  9.850000n 0.9  9.875000n 0.9  9.975000n 0.9  10.000000n 0.9  10.100000n 0.9  10.125000n 0.9  10.225000n 0.9  10.250000n 0.9  10.350000n 0.9  10.375000n 0.9  10.475000n 0.9  10.500000n 0.9  10.600000n 0.9  10.625000n 0.9  10.725000n 0.9  10.750000n 0.9  10.850000n 0.9  10.875000n 0.9  10.975000n 0.9  11.000000n 0.9  11.100000n 0.9  11.125000n 0.9  11.225000n 0.9  11.250000n 0.0  11.350000n 0.0  11.375000n 0.0  11.475000n 0.0  11.500000n 0.0  11.600000n 0.0  11.625000n 0.0  11.725000n 0.0  11.750000n 0.0  11.850000n 0.0  11.875000n 0.0  11.975000n 0.0  12.000000n 0.0  12.100000n 0.0  12.125000n 0.0  12.225000n 0.0  12.250000n 0.0  12.350000n 0.0  12.375000n 0.0  12.475000n 0.0  12.500000n 0.0  12.600000n 0.0  12.625000n 0.0  12.725000n 0.0  12.750000n 0.0  12.850000n 0.0  12.875000n 0.0  12.975000n 0.0  13.000000n 0.0  13.100000n 0.0  13.125000n 0.0  13.225000n 0.0  13.250000n 0.0  13.350000n 0.0  13.375000n 0.0  13.475000n 0.0  13.500000n 0.0  13.600000n 0.0  13.625000n 0.0  13.725000n 0.0  13.750000n 0.0  13.850000n 0.0  13.875000n 0.0  13.975000n 0.0  14.000000n 0.0  14.100000n 0.0  14.125000n 0.0  14.225000n 0.0  14.250000n 0.0  14.350000n 0.0  14.375000n 0.0  14.475000n 0.0  14.500000n 0.0  14.600000n 0.0  14.625000n 0.0  14.725000n 0.0  14.750000n 0.0  14.850000n 0.0  14.875000n 0.0  14.975000n 0.0  15.000000n 0.0  15.100000n 0.0  15.125000n 0.0  15.225000n 0.0  15.250000n 0.0  15.350000n 0.0  15.375000n 0.0  15.475000n 0.0  15.500000n 0.0  15.600000n 0.0  15.625000n 0.0  15.725000n 0.0  15.750000n 0.9  15.850000n 0.9  15.875000n 0.9  15.975000n 0.9  16.000000n 0.9  16.100000n 0.9  16.125000n 0.9  16.225000n 0.9  16.250000n 0.9  16.350000n 0.9  16.375000n 0.9  16.475000n 0.9  16.500000n 0.9  16.600000n 0.9  16.625000n 0.9  16.725000n 0.9  16.750000n 0.9  16.850000n 0.9  16.875000n 0.9  16.975000n 0.9  17.000000n 0.9  17.100000n 0.9  17.125000n 0.9  17.225000n 0.9  17.250000n 0.9  17.350000n 0.9  17.375000n 0.9  17.475000n 0.9  17.500000n 0.9  17.600000n 0.9  17.625000n 0.9  17.725000n 0.9  17.750000n 0.9  17.850000n 0.9  17.875000n 0.9  17.975000n 0.9  18.000000n 0.0  18.100000n 0.0  18.125000n 0.0  18.225000n 0.0  18.250000n 0.0  18.350000n 0.0  18.375000n 0.0  18.475000n 0.0  18.500000n 0.0  18.600000n 0.0  18.625000n 0.0  18.725000n 0.0  18.750000n 0.0  18.850000n 0.0  18.875000n 0.0  18.975000n 0.0  19.000000n 0.0  19.100000n 0.0  19.125000n 0.0  19.225000n 0.0  19.250000n 0.0  19.350000n 0.0  19.375000n 0.0  19.475000n 0.0  19.500000n 0.0  19.600000n 0.0  19.625000n 0.0  19.725000n 0.0  19.750000n 0.0  19.850000n 0.0  19.875000n 0.0  19.975000n 0.0  20.000000n 0.0  20.100000n 0.0  20.125000n 0.0  20.225000n 0.0  20.250000n 0.0  20.350000n 0.0  20.375000n 0.0  20.475000n 0.0  20.500000n 0.0  20.600000n 0.0  20.625000n 0.0  20.725000n 0.0  20.750000n 0.0  20.850000n 0.0  20.875000n 0.0  20.975000n 0.0  21.000000n 0.0  21.100000n 0.0  21.125000n 0.0  21.225000n 0.0  21.250000n 0.0  21.350000n 0.0  21.375000n 0.0  21.475000n 0.0  21.500000n 0.0  21.600000n 0.0  21.625000n 0.0  21.725000n 0.0  21.750000n 0.0  21.850000n 0.0  21.875000n 0.0  21.975000n 0.0  22.000000n 0.0  22.100000n 0.0  22.125000n 0.0  22.225000n 0.0  22.250000n 0.0  22.350000n 0.0  22.375000n 0.0  22.475000n 0.0  22.500000n 0.9  22.600000n 0.9  22.625000n 0.9  22.725000n 0.9  22.750000n 0.9  22.850000n 0.9  22.875000n 0.9  22.975000n 0.9  23.000000n 0.9  23.100000n 0.9  23.125000n 0.9  23.225000n 0.9  23.250000n 0.9  23.350000n 0.9  23.375000n 0.9  23.475000n 0.9  23.500000n 0.9  23.600000n 0.9  23.625000n 0.9  23.725000n 0.9  23.750000n 0.9  23.850000n 0.9  23.875000n 0.9  23.975000n 0.9  24.000000n 0.9  24.100000n 0.9  24.125000n 0.9  24.225000n 0.9  24.250000n 0.9  24.350000n 0.9  24.375000n 0.9  24.475000n 0.9  24.500000n 0.9  24.600000n 0.9  24.625000n 0.9  24.725000n 0.9  24.750000n 0.0  24.850000n 0.0  24.875000n 0.0  24.975000n 0.0  25.000000n 0.0  25.100000n 0.0  25.125000n 0.0  25.225000n 0.0  25.250000n 0.0  25.350000n 0.0  25.375000n 0.0  25.475000n 0.0  25.500000n 0.0  25.600000n 0.0  25.625000n 0.0  25.725000n 0.0  25.750000n 0.0  25.850000n 0.0  25.875000n 0.0  25.975000n 0.0  26.000000n 0.0  26.100000n 0.0  26.125000n 0.0  26.225000n 0.0  26.250000n 0.0  26.350000n 0.0  26.375000n 0.0  26.475000n 0.0  26.500000n 0.0  26.600000n 0.0  26.625000n 0.0  26.725000n 0.0  26.750000n 0.0  26.850000n 0.0  26.875000n 0.0  26.975000n 0.0  27.000000n 0.0  27.100000n 0.0  27.125000n 0.0  27.225000n 0.0  27.250000n 0.0  27.350000n 0.0  27.375000n 0.0  27.475000n 0.0  27.500000n 0.0  27.600000n 0.0  27.625000n 0.0  27.725000n 0.0  27.750000n 0.0  27.850000n 0.0  27.875000n 0.0  27.975000n 0.0  28.000000n 0.0  28.100000n 0.0  28.125000n 0.0  28.225000n 0.0  28.250000n 0.0  28.350000n 0.0  28.375000n 0.0  28.475000n 0.0  28.500000n 0.0  28.600000n 0.0  28.625000n 0.0  28.725000n 0.0  28.750000n 0.0  28.850000n 0.0  28.875000n 0.0  28.975000n 0.0  29.000000n 0.0  29.100000n 0.0  29.125000n 0.0  29.225000n 0.0  29.250000n 0.9  29.350000n 0.9  29.375000n 0.9  29.475000n 0.9  29.500000n 0.9  29.600000n 0.9  29.625000n 0.9  29.725000n 0.9  29.750000n 0.9  29.850000n 0.9  29.875000n 0.9  29.975000n 0.9  30.000000n 0.9  30.100000n 0.9  30.125000n 0.9  30.225000n 0.9  30.250000n 0.9 )
V_W00<0> W00<0> 0 PWL(0.000000n 0.0  0.100000n 0.0  0.125000n 0.0  0.225000n 0.0  0.250000n 0.0  0.350000n 0.0  0.375000n 0.0  0.475000n 0.0  0.500000n 0.0  0.600000n 0.0  0.625000n 0.0  0.725000n 0.0  0.750000n 0.0  0.850000n 0.0  0.875000n 0.0  0.975000n 0.0  1.000000n 0.0  1.100000n 0.0  1.125000n 0.9  1.225000n 0.9  1.250000n 0.9  1.350000n 0.9  1.375000n 0.9  1.475000n 0.9  1.500000n 0.9  1.600000n 0.9  1.625000n 0.9  1.725000n 0.9  1.750000n 0.9  1.850000n 0.9  1.875000n 0.9  1.975000n 0.9  2.000000n 0.9  2.100000n 0.9  2.125000n 0.9  2.225000n 0.9  2.250000n 0.9  2.350000n 0.9  2.375000n 0.9  2.475000n 0.9  2.500000n 0.9  2.600000n 0.9  2.625000n 0.9  2.725000n 0.9  2.750000n 0.9  2.850000n 0.9  2.875000n 0.9  2.975000n 0.9  3.000000n 0.9  3.100000n 0.9  3.125000n 0.9  3.225000n 0.9  3.250000n 0.9  3.350000n 0.9  3.375000n 0.9  3.475000n 0.9  3.500000n 0.9  3.600000n 0.9  3.625000n 0.9  3.725000n 0.9  3.750000n 0.9  3.850000n 0.9  3.875000n 0.9  3.975000n 0.9  4.000000n 0.9  4.100000n 0.9  4.125000n 0.9  4.225000n 0.9  4.250000n 0.9  4.350000n 0.9  4.375000n 0.9  4.475000n 0.9  4.500000n 0.9  4.600000n 0.9  4.625000n 0.9  4.725000n 0.9  4.750000n 0.9  4.850000n 0.9  4.875000n 0.9  4.975000n 0.9  5.000000n 0.9  5.100000n 0.9  5.125000n 0.9  5.225000n 0.9  5.250000n 0.9  5.350000n 0.9  5.375000n 0.9  5.475000n 0.9  5.500000n 0.9  5.600000n 0.9  5.625000n 0.0  5.725000n 0.0  5.750000n 0.0  5.850000n 0.0  5.875000n 0.0  5.975000n 0.0  6.000000n 0.0  6.100000n 0.0  6.125000n 0.0  6.225000n 0.0  6.250000n 0.0  6.350000n 0.0  6.375000n 0.0  6.475000n 0.0  6.500000n 0.0  6.600000n 0.0  6.625000n 0.0  6.725000n 0.0  6.750000n 0.0  6.850000n 0.0  6.875000n 0.0  6.975000n 0.0  7.000000n 0.0  7.100000n 0.0  7.125000n 0.0  7.225000n 0.0  7.250000n 0.0  7.350000n 0.0  7.375000n 0.0  7.475000n 0.0  7.500000n 0.0  7.600000n 0.0  7.625000n 0.0  7.725000n 0.0  7.750000n 0.0  7.850000n 0.0  7.875000n 0.9  7.975000n 0.9  8.000000n 0.9  8.100000n 0.9  8.125000n 0.9  8.225000n 0.9  8.250000n 0.9  8.350000n 0.9  8.375000n 0.9  8.475000n 0.9  8.500000n 0.9  8.600000n 0.9  8.625000n 0.9  8.725000n 0.9  8.750000n 0.9  8.850000n 0.9  8.875000n 0.9  8.975000n 0.9  9.000000n 0.9  9.100000n 0.9  9.125000n 0.9  9.225000n 0.9  9.250000n 0.9  9.350000n 0.9  9.375000n 0.9  9.475000n 0.9  9.500000n 0.9  9.600000n 0.9  9.625000n 0.9  9.725000n 0.9  9.750000n 0.9  9.850000n 0.9  9.875000n 0.9  9.975000n 0.9  10.000000n 0.9  10.100000n 0.9  10.125000n 0.9  10.225000n 0.9  10.250000n 0.9  10.350000n 0.9  10.375000n 0.9  10.475000n 0.9  10.500000n 0.9  10.600000n 0.9  10.625000n 0.9  10.725000n 0.9  10.750000n 0.9  10.850000n 0.9  10.875000n 0.9  10.975000n 0.9  11.000000n 0.9  11.100000n 0.9  11.125000n 0.9  11.225000n 0.9  11.250000n 0.9  11.350000n 0.9  11.375000n 0.9  11.475000n 0.9  11.500000n 0.9  11.600000n 0.9  11.625000n 0.9  11.725000n 0.9  11.750000n 0.9  11.850000n 0.9  11.875000n 0.9  11.975000n 0.9  12.000000n 0.9  12.100000n 0.9  12.125000n 0.9  12.225000n 0.9  12.250000n 0.9  12.350000n 0.9  12.375000n 0.0  12.475000n 0.0  12.500000n 0.0  12.600000n 0.0  12.625000n 0.0  12.725000n 0.0  12.750000n 0.0  12.850000n 0.0  12.875000n 0.0  12.975000n 0.0  13.000000n 0.0  13.100000n 0.0  13.125000n 0.0  13.225000n 0.0  13.250000n 0.0  13.350000n 0.0  13.375000n 0.0  13.475000n 0.0  13.500000n 0.0  13.600000n 0.0  13.625000n 0.0  13.725000n 0.0  13.750000n 0.0  13.850000n 0.0  13.875000n 0.0  13.975000n 0.0  14.000000n 0.0  14.100000n 0.0  14.125000n 0.0  14.225000n 0.0  14.250000n 0.0  14.350000n 0.0  14.375000n 0.0  14.475000n 0.0  14.500000n 0.0  14.600000n 0.0  14.625000n 0.9  14.725000n 0.9  14.750000n 0.9  14.850000n 0.9  14.875000n 0.9  14.975000n 0.9  15.000000n 0.9  15.100000n 0.9  15.125000n 0.9  15.225000n 0.9  15.250000n 0.9  15.350000n 0.9  15.375000n 0.9  15.475000n 0.9  15.500000n 0.9  15.600000n 0.9  15.625000n 0.9  15.725000n 0.9  15.750000n 0.9  15.850000n 0.9  15.875000n 0.9  15.975000n 0.9  16.000000n 0.9  16.100000n 0.9  16.125000n 0.9  16.225000n 0.9  16.250000n 0.9  16.350000n 0.9  16.375000n 0.9  16.475000n 0.9  16.500000n 0.9  16.600000n 0.9  16.625000n 0.9  16.725000n 0.9  16.750000n 0.9  16.850000n 0.9  16.875000n 0.9  16.975000n 0.9  17.000000n 0.9  17.100000n 0.9  17.125000n 0.9  17.225000n 0.9  17.250000n 0.9  17.350000n 0.9  17.375000n 0.9  17.475000n 0.9  17.500000n 0.9  17.600000n 0.9  17.625000n 0.9  17.725000n 0.9  17.750000n 0.9  17.850000n 0.9  17.875000n 0.9  17.975000n 0.9  18.000000n 0.9  18.100000n 0.9  18.125000n 0.9  18.225000n 0.9  18.250000n 0.9  18.350000n 0.9  18.375000n 0.9  18.475000n 0.9  18.500000n 0.9  18.600000n 0.9  18.625000n 0.9  18.725000n 0.9  18.750000n 0.9  18.850000n 0.9  18.875000n 0.9  18.975000n 0.9  19.000000n 0.9  19.100000n 0.9  19.125000n 0.0  19.225000n 0.0  19.250000n 0.0  19.350000n 0.0  19.375000n 0.0  19.475000n 0.0  19.500000n 0.0  19.600000n 0.0  19.625000n 0.0  19.725000n 0.0  19.750000n 0.0  19.850000n 0.0  19.875000n 0.0  19.975000n 0.0  20.000000n 0.0  20.100000n 0.0  20.125000n 0.0  20.225000n 0.0  20.250000n 0.0  20.350000n 0.0  20.375000n 0.0  20.475000n 0.0  20.500000n 0.0  20.600000n 0.0  20.625000n 0.0  20.725000n 0.0  20.750000n 0.0  20.850000n 0.0  20.875000n 0.0  20.975000n 0.0  21.000000n 0.0  21.100000n 0.0  21.125000n 0.0  21.225000n 0.0  21.250000n 0.0  21.350000n 0.0  21.375000n 0.9  21.475000n 0.9  21.500000n 0.9  21.600000n 0.9  21.625000n 0.9  21.725000n 0.9  21.750000n 0.9  21.850000n 0.9  21.875000n 0.9  21.975000n 0.9  22.000000n 0.9  22.100000n 0.9  22.125000n 0.9  22.225000n 0.9  22.250000n 0.9  22.350000n 0.9  22.375000n 0.9  22.475000n 0.9  22.500000n 0.9  22.600000n 0.9  22.625000n 0.9  22.725000n 0.9  22.750000n 0.9  22.850000n 0.9  22.875000n 0.9  22.975000n 0.9  23.000000n 0.9  23.100000n 0.9  23.125000n 0.9  23.225000n 0.9  23.250000n 0.9  23.350000n 0.9  23.375000n 0.9  23.475000n 0.9  23.500000n 0.9  23.600000n 0.9  23.625000n 0.9  23.725000n 0.9  23.750000n 0.9  23.850000n 0.9  23.875000n 0.9  23.975000n 0.9  24.000000n 0.9  24.100000n 0.9  24.125000n 0.9  24.225000n 0.9  24.250000n 0.9  24.350000n 0.9  24.375000n 0.9  24.475000n 0.9  24.500000n 0.9  24.600000n 0.9  24.625000n 0.9  24.725000n 0.9  24.750000n 0.9  24.850000n 0.9  24.875000n 0.9  24.975000n 0.9  25.000000n 0.9  25.100000n 0.9  25.125000n 0.9  25.225000n 0.9  25.250000n 0.9  25.350000n 0.9  25.375000n 0.9  25.475000n 0.9  25.500000n 0.9  25.600000n 0.9  25.625000n 0.9  25.725000n 0.9  25.750000n 0.9  25.850000n 0.9  25.875000n 0.0  25.975000n 0.0  26.000000n 0.0  26.100000n 0.0  26.125000n 0.0  26.225000n 0.0  26.250000n 0.0  26.350000n 0.0  26.375000n 0.0  26.475000n 0.0  26.500000n 0.0  26.600000n 0.0  26.625000n 0.0  26.725000n 0.0  26.750000n 0.0  26.850000n 0.0  26.875000n 0.0  26.975000n 0.0  27.000000n 0.0  27.100000n 0.0  27.125000n 0.0  27.225000n 0.0  27.250000n 0.0  27.350000n 0.0  27.375000n 0.0  27.475000n 0.0  27.500000n 0.0  27.600000n 0.0  27.625000n 0.0  27.725000n 0.0  27.750000n 0.0  27.850000n 0.0  27.875000n 0.0  27.975000n 0.0  28.000000n 0.0  28.100000n 0.0  28.125000n 0.9  28.225000n 0.9  28.250000n 0.9  28.350000n 0.9  28.375000n 0.9  28.475000n 0.9  28.500000n 0.9  28.600000n 0.9  28.625000n 0.9  28.725000n 0.9  28.750000n 0.9  28.850000n 0.9  28.875000n 0.9  28.975000n 0.9  29.000000n 0.9  29.100000n 0.9  29.125000n 0.9  29.225000n 0.9  29.250000n 0.9  29.350000n 0.9  29.375000n 0.9  29.475000n 0.9  29.500000n 0.9  29.600000n 0.9  29.625000n 0.9  29.725000n 0.9  29.750000n 0.9  29.850000n 0.9  29.875000n 0.9  29.975000n 0.9  30.000000n 0.9  30.100000n 0.9  30.125000n 0.9  30.225000n 0.9  30.250000n 0.9 )
V_W01<1> W01<1> 0 PWL(0.000000n 0.0  0.100000n 0.0  0.125000n 0.0  0.225000n 0.0  0.250000n 0.0  0.350000n 0.0  0.375000n 0.0  0.475000n 0.0  0.500000n 0.0  0.600000n 0.0  0.625000n 0.0  0.725000n 0.0  0.750000n 0.9  0.850000n 0.9  0.875000n 0.9  0.975000n 0.9  1.000000n 0.9  1.100000n 0.9  1.125000n 0.9  1.225000n 0.9  1.250000n 0.9  1.350000n 0.9  1.375000n 0.9  1.475000n 0.9  1.500000n 0.0  1.600000n 0.0  1.625000n 0.0  1.725000n 0.0  1.750000n 0.0  1.850000n 0.0  1.875000n 0.0  1.975000n 0.0  2.000000n 0.0  2.100000n 0.0  2.125000n 0.0  2.225000n 0.0  2.250000n 0.0  2.350000n 0.0  2.375000n 0.0  2.475000n 0.0  2.500000n 0.0  2.600000n 0.0  2.625000n 0.0  2.725000n 0.0  2.750000n 0.0  2.850000n 0.0  2.875000n 0.0  2.975000n 0.0  3.000000n 0.9  3.100000n 0.9  3.125000n 0.9  3.225000n 0.9  3.250000n 0.9  3.350000n 0.9  3.375000n 0.9  3.475000n 0.9  3.500000n 0.9  3.600000n 0.9  3.625000n 0.9  3.725000n 0.9  3.750000n 0.0  3.850000n 0.0  3.875000n 0.0  3.975000n 0.0  4.000000n 0.0  4.100000n 0.0  4.125000n 0.0  4.225000n 0.0  4.250000n 0.0  4.350000n 0.0  4.375000n 0.0  4.475000n 0.0  4.500000n 0.0  4.600000n 0.0  4.625000n 0.0  4.725000n 0.0  4.750000n 0.0  4.850000n 0.0  4.875000n 0.0  4.975000n 0.0  5.000000n 0.0  5.100000n 0.0  5.125000n 0.0  5.225000n 0.0  5.250000n 0.9  5.350000n 0.9  5.375000n 0.9  5.475000n 0.9  5.500000n 0.9  5.600000n 0.9  5.625000n 0.9  5.725000n 0.9  5.750000n 0.9  5.850000n 0.9  5.875000n 0.9  5.975000n 0.9  6.000000n 0.0  6.100000n 0.0  6.125000n 0.0  6.225000n 0.0  6.250000n 0.0  6.350000n 0.0  6.375000n 0.0  6.475000n 0.0  6.500000n 0.0  6.600000n 0.0  6.625000n 0.0  6.725000n 0.0  6.750000n 0.0  6.850000n 0.0  6.875000n 0.0  6.975000n 0.0  7.000000n 0.0  7.100000n 0.0  7.125000n 0.0  7.225000n 0.0  7.250000n 0.0  7.350000n 0.0  7.375000n 0.0  7.475000n 0.0  7.500000n 0.9  7.600000n 0.9  7.625000n 0.9  7.725000n 0.9  7.750000n 0.9  7.850000n 0.9  7.875000n 0.9  7.975000n 0.9  8.000000n 0.9  8.100000n 0.9  8.125000n 0.9  8.225000n 0.9  8.250000n 0.0  8.350000n 0.0  8.375000n 0.0  8.475000n 0.0  8.500000n 0.0  8.600000n 0.0  8.625000n 0.0  8.725000n 0.0  8.750000n 0.0  8.850000n 0.0  8.875000n 0.0  8.975000n 0.0  9.000000n 0.0  9.100000n 0.0  9.125000n 0.0  9.225000n 0.0  9.250000n 0.0  9.350000n 0.0  9.375000n 0.0  9.475000n 0.0  9.500000n 0.0  9.600000n 0.0  9.625000n 0.0  9.725000n 0.0  9.750000n 0.9  9.850000n 0.9  9.875000n 0.9  9.975000n 0.9  10.000000n 0.9  10.100000n 0.9  10.125000n 0.9  10.225000n 0.9  10.250000n 0.9  10.350000n 0.9  10.375000n 0.9  10.475000n 0.9  10.500000n 0.0  10.600000n 0.0  10.625000n 0.0  10.725000n 0.0  10.750000n 0.0  10.850000n 0.0  10.875000n 0.0  10.975000n 0.0  11.000000n 0.0  11.100000n 0.0  11.125000n 0.0  11.225000n 0.0  11.250000n 0.0  11.350000n 0.0  11.375000n 0.0  11.475000n 0.0  11.500000n 0.0  11.600000n 0.0  11.625000n 0.0  11.725000n 0.0  11.750000n 0.0  11.850000n 0.0  11.875000n 0.0  11.975000n 0.0  12.000000n 0.9  12.100000n 0.9  12.125000n 0.9  12.225000n 0.9  12.250000n 0.9  12.350000n 0.9  12.375000n 0.9  12.475000n 0.9  12.500000n 0.9  12.600000n 0.9  12.625000n 0.9  12.725000n 0.9  12.750000n 0.0  12.850000n 0.0  12.875000n 0.0  12.975000n 0.0  13.000000n 0.0  13.100000n 0.0  13.125000n 0.0  13.225000n 0.0  13.250000n 0.0  13.350000n 0.0  13.375000n 0.0  13.475000n 0.0  13.500000n 0.0  13.600000n 0.0  13.625000n 0.0  13.725000n 0.0  13.750000n 0.0  13.850000n 0.0  13.875000n 0.0  13.975000n 0.0  14.000000n 0.0  14.100000n 0.0  14.125000n 0.0  14.225000n 0.0  14.250000n 0.9  14.350000n 0.9  14.375000n 0.9  14.475000n 0.9  14.500000n 0.9  14.600000n 0.9  14.625000n 0.9  14.725000n 0.9  14.750000n 0.9  14.850000n 0.9  14.875000n 0.9  14.975000n 0.9  15.000000n 0.0  15.100000n 0.0  15.125000n 0.0  15.225000n 0.0  15.250000n 0.0  15.350000n 0.0  15.375000n 0.0  15.475000n 0.0  15.500000n 0.0  15.600000n 0.0  15.625000n 0.0  15.725000n 0.0  15.750000n 0.0  15.850000n 0.0  15.875000n 0.0  15.975000n 0.0  16.000000n 0.0  16.100000n 0.0  16.125000n 0.0  16.225000n 0.0  16.250000n 0.0  16.350000n 0.0  16.375000n 0.0  16.475000n 0.0  16.500000n 0.9  16.600000n 0.9  16.625000n 0.9  16.725000n 0.9  16.750000n 0.9  16.850000n 0.9  16.875000n 0.9  16.975000n 0.9  17.000000n 0.9  17.100000n 0.9  17.125000n 0.9  17.225000n 0.9  17.250000n 0.0  17.350000n 0.0  17.375000n 0.0  17.475000n 0.0  17.500000n 0.0  17.600000n 0.0  17.625000n 0.0  17.725000n 0.0  17.750000n 0.0  17.850000n 0.0  17.875000n 0.0  17.975000n 0.0  18.000000n 0.0  18.100000n 0.0  18.125000n 0.0  18.225000n 0.0  18.250000n 0.0  18.350000n 0.0  18.375000n 0.0  18.475000n 0.0  18.500000n 0.0  18.600000n 0.0  18.625000n 0.0  18.725000n 0.0  18.750000n 0.9  18.850000n 0.9  18.875000n 0.9  18.975000n 0.9  19.000000n 0.9  19.100000n 0.9  19.125000n 0.9  19.225000n 0.9  19.250000n 0.9  19.350000n 0.9  19.375000n 0.9  19.475000n 0.9  19.500000n 0.0  19.600000n 0.0  19.625000n 0.0  19.725000n 0.0  19.750000n 0.0  19.850000n 0.0  19.875000n 0.0  19.975000n 0.0  20.000000n 0.0  20.100000n 0.0  20.125000n 0.0  20.225000n 0.0  20.250000n 0.0  20.350000n 0.0  20.375000n 0.0  20.475000n 0.0  20.500000n 0.0  20.600000n 0.0  20.625000n 0.0  20.725000n 0.0  20.750000n 0.0  20.850000n 0.0  20.875000n 0.0  20.975000n 0.0  21.000000n 0.9  21.100000n 0.9  21.125000n 0.9  21.225000n 0.9  21.250000n 0.9  21.350000n 0.9  21.375000n 0.9  21.475000n 0.9  21.500000n 0.9  21.600000n 0.9  21.625000n 0.9  21.725000n 0.9  21.750000n 0.0  21.850000n 0.0  21.875000n 0.0  21.975000n 0.0  22.000000n 0.0  22.100000n 0.0  22.125000n 0.0  22.225000n 0.0  22.250000n 0.0  22.350000n 0.0  22.375000n 0.0  22.475000n 0.0  22.500000n 0.0  22.600000n 0.0  22.625000n 0.0  22.725000n 0.0  22.750000n 0.0  22.850000n 0.0  22.875000n 0.0  22.975000n 0.0  23.000000n 0.0  23.100000n 0.0  23.125000n 0.0  23.225000n 0.0  23.250000n 0.9  23.350000n 0.9  23.375000n 0.9  23.475000n 0.9  23.500000n 0.9  23.600000n 0.9  23.625000n 0.9  23.725000n 0.9  23.750000n 0.9  23.850000n 0.9  23.875000n 0.9  23.975000n 0.9  24.000000n 0.0  24.100000n 0.0  24.125000n 0.0  24.225000n 0.0  24.250000n 0.0  24.350000n 0.0  24.375000n 0.0  24.475000n 0.0  24.500000n 0.0  24.600000n 0.0  24.625000n 0.0  24.725000n 0.0  24.750000n 0.0  24.850000n 0.0  24.875000n 0.0  24.975000n 0.0  25.000000n 0.0  25.100000n 0.0  25.125000n 0.0  25.225000n 0.0  25.250000n 0.0  25.350000n 0.0  25.375000n 0.0  25.475000n 0.0  25.500000n 0.9  25.600000n 0.9  25.625000n 0.9  25.725000n 0.9  25.750000n 0.9  25.850000n 0.9  25.875000n 0.9  25.975000n 0.9  26.000000n 0.9  26.100000n 0.9  26.125000n 0.9  26.225000n 0.9  26.250000n 0.0  26.350000n 0.0  26.375000n 0.0  26.475000n 0.0  26.500000n 0.0  26.600000n 0.0  26.625000n 0.0  26.725000n 0.0  26.750000n 0.0  26.850000n 0.0  26.875000n 0.0  26.975000n 0.0  27.000000n 0.0  27.100000n 0.0  27.125000n 0.0  27.225000n 0.0  27.250000n 0.0  27.350000n 0.0  27.375000n 0.0  27.475000n 0.0  27.500000n 0.0  27.600000n 0.0  27.625000n 0.0  27.725000n 0.0  27.750000n 0.9  27.850000n 0.9  27.875000n 0.9  27.975000n 0.9  28.000000n 0.9  28.100000n 0.9  28.125000n 0.9  28.225000n 0.9  28.250000n 0.9  28.350000n 0.9  28.375000n 0.9  28.475000n 0.9  28.500000n 0.0  28.600000n 0.0  28.625000n 0.0  28.725000n 0.0  28.750000n 0.0  28.850000n 0.0  28.875000n 0.0  28.975000n 0.0  29.000000n 0.0  29.100000n 0.0  29.125000n 0.0  29.225000n 0.0  29.250000n 0.0  29.350000n 0.0  29.375000n 0.0  29.475000n 0.0  29.500000n 0.0  29.600000n 0.0  29.625000n 0.0  29.725000n 0.0  29.750000n 0.0  29.850000n 0.0  29.875000n 0.0  29.975000n 0.0  30.000000n 0.9  30.100000n 0.9  30.125000n 0.9  30.225000n 0.9  30.250000n 0.9 )
V_W01<0> W01<0> 0 PWL(0.000000n 0.0  0.100000n 0.0  0.125000n 0.0  0.225000n 0.0  0.250000n 0.0  0.350000n 0.0  0.375000n 0.9  0.475000n 0.9  0.500000n 0.9  0.600000n 0.9  0.625000n 0.9  0.725000n 0.9  0.750000n 0.9  0.850000n 0.9  0.875000n 0.9  0.975000n 0.9  1.000000n 0.9  1.100000n 0.9  1.125000n 0.9  1.225000n 0.9  1.250000n 0.9  1.350000n 0.9  1.375000n 0.9  1.475000n 0.9  1.500000n 0.9  1.600000n 0.9  1.625000n 0.9  1.725000n 0.9  1.750000n 0.9  1.850000n 0.9  1.875000n 0.0  1.975000n 0.0  2.000000n 0.0  2.100000n 0.0  2.125000n 0.0  2.225000n 0.0  2.250000n 0.0  2.350000n 0.0  2.375000n 0.0  2.475000n 0.0  2.500000n 0.0  2.600000n 0.0  2.625000n 0.9  2.725000n 0.9  2.750000n 0.9  2.850000n 0.9  2.875000n 0.9  2.975000n 0.9  3.000000n 0.9  3.100000n 0.9  3.125000n 0.9  3.225000n 0.9  3.250000n 0.9  3.350000n 0.9  3.375000n 0.9  3.475000n 0.9  3.500000n 0.9  3.600000n 0.9  3.625000n 0.9  3.725000n 0.9  3.750000n 0.9  3.850000n 0.9  3.875000n 0.9  3.975000n 0.9  4.000000n 0.9  4.100000n 0.9  4.125000n 0.0  4.225000n 0.0  4.250000n 0.0  4.350000n 0.0  4.375000n 0.0  4.475000n 0.0  4.500000n 0.0  4.600000n 0.0  4.625000n 0.0  4.725000n 0.0  4.750000n 0.0  4.850000n 0.0  4.875000n 0.9  4.975000n 0.9  5.000000n 0.9  5.100000n 0.9  5.125000n 0.9  5.225000n 0.9  5.250000n 0.9  5.350000n 0.9  5.375000n 0.9  5.475000n 0.9  5.500000n 0.9  5.600000n 0.9  5.625000n 0.9  5.725000n 0.9  5.750000n 0.9  5.850000n 0.9  5.875000n 0.9  5.975000n 0.9  6.000000n 0.9  6.100000n 0.9  6.125000n 0.9  6.225000n 0.9  6.250000n 0.9  6.350000n 0.9  6.375000n 0.0  6.475000n 0.0  6.500000n 0.0  6.600000n 0.0  6.625000n 0.0  6.725000n 0.0  6.750000n 0.0  6.850000n 0.0  6.875000n 0.0  6.975000n 0.0  7.000000n 0.0  7.100000n 0.0  7.125000n 0.9  7.225000n 0.9  7.250000n 0.9  7.350000n 0.9  7.375000n 0.9  7.475000n 0.9  7.500000n 0.9  7.600000n 0.9  7.625000n 0.9  7.725000n 0.9  7.750000n 0.9  7.850000n 0.9  7.875000n 0.9  7.975000n 0.9  8.000000n 0.9  8.100000n 0.9  8.125000n 0.9  8.225000n 0.9  8.250000n 0.9  8.350000n 0.9  8.375000n 0.9  8.475000n 0.9  8.500000n 0.9  8.600000n 0.9  8.625000n 0.0  8.725000n 0.0  8.750000n 0.0  8.850000n 0.0  8.875000n 0.0  8.975000n 0.0  9.000000n 0.0  9.100000n 0.0  9.125000n 0.0  9.225000n 0.0  9.250000n 0.0  9.350000n 0.0  9.375000n 0.9  9.475000n 0.9  9.500000n 0.9  9.600000n 0.9  9.625000n 0.9  9.725000n 0.9  9.750000n 0.9  9.850000n 0.9  9.875000n 0.9  9.975000n 0.9  10.000000n 0.9  10.100000n 0.9  10.125000n 0.9  10.225000n 0.9  10.250000n 0.9  10.350000n 0.9  10.375000n 0.9  10.475000n 0.9  10.500000n 0.9  10.600000n 0.9  10.625000n 0.9  10.725000n 0.9  10.750000n 0.9  10.850000n 0.9  10.875000n 0.0  10.975000n 0.0  11.000000n 0.0  11.100000n 0.0  11.125000n 0.0  11.225000n 0.0  11.250000n 0.0  11.350000n 0.0  11.375000n 0.0  11.475000n 0.0  11.500000n 0.0  11.600000n 0.0  11.625000n 0.9  11.725000n 0.9  11.750000n 0.9  11.850000n 0.9  11.875000n 0.9  11.975000n 0.9  12.000000n 0.9  12.100000n 0.9  12.125000n 0.9  12.225000n 0.9  12.250000n 0.9  12.350000n 0.9  12.375000n 0.9  12.475000n 0.9  12.500000n 0.9  12.600000n 0.9  12.625000n 0.9  12.725000n 0.9  12.750000n 0.9  12.850000n 0.9  12.875000n 0.9  12.975000n 0.9  13.000000n 0.9  13.100000n 0.9  13.125000n 0.0  13.225000n 0.0  13.250000n 0.0  13.350000n 0.0  13.375000n 0.0  13.475000n 0.0  13.500000n 0.0  13.600000n 0.0  13.625000n 0.0  13.725000n 0.0  13.750000n 0.0  13.850000n 0.0  13.875000n 0.9  13.975000n 0.9  14.000000n 0.9  14.100000n 0.9  14.125000n 0.9  14.225000n 0.9  14.250000n 0.9  14.350000n 0.9  14.375000n 0.9  14.475000n 0.9  14.500000n 0.9  14.600000n 0.9  14.625000n 0.9  14.725000n 0.9  14.750000n 0.9  14.850000n 0.9  14.875000n 0.9  14.975000n 0.9  15.000000n 0.9  15.100000n 0.9  15.125000n 0.9  15.225000n 0.9  15.250000n 0.9  15.350000n 0.9  15.375000n 0.0  15.475000n 0.0  15.500000n 0.0  15.600000n 0.0  15.625000n 0.0  15.725000n 0.0  15.750000n 0.0  15.850000n 0.0  15.875000n 0.0  15.975000n 0.0  16.000000n 0.0  16.100000n 0.0  16.125000n 0.9  16.225000n 0.9  16.250000n 0.9  16.350000n 0.9  16.375000n 0.9  16.475000n 0.9  16.500000n 0.9  16.600000n 0.9  16.625000n 0.9  16.725000n 0.9  16.750000n 0.9  16.850000n 0.9  16.875000n 0.9  16.975000n 0.9  17.000000n 0.9  17.100000n 0.9  17.125000n 0.9  17.225000n 0.9  17.250000n 0.9  17.350000n 0.9  17.375000n 0.9  17.475000n 0.9  17.500000n 0.9  17.600000n 0.9  17.625000n 0.0  17.725000n 0.0  17.750000n 0.0  17.850000n 0.0  17.875000n 0.0  17.975000n 0.0  18.000000n 0.0  18.100000n 0.0  18.125000n 0.0  18.225000n 0.0  18.250000n 0.0  18.350000n 0.0  18.375000n 0.9  18.475000n 0.9  18.500000n 0.9  18.600000n 0.9  18.625000n 0.9  18.725000n 0.9  18.750000n 0.9  18.850000n 0.9  18.875000n 0.9  18.975000n 0.9  19.000000n 0.9  19.100000n 0.9  19.125000n 0.9  19.225000n 0.9  19.250000n 0.9  19.350000n 0.9  19.375000n 0.9  19.475000n 0.9  19.500000n 0.9  19.600000n 0.9  19.625000n 0.9  19.725000n 0.9  19.750000n 0.9  19.850000n 0.9  19.875000n 0.0  19.975000n 0.0  20.000000n 0.0  20.100000n 0.0  20.125000n 0.0  20.225000n 0.0  20.250000n 0.0  20.350000n 0.0  20.375000n 0.0  20.475000n 0.0  20.500000n 0.0  20.600000n 0.0  20.625000n 0.9  20.725000n 0.9  20.750000n 0.9  20.850000n 0.9  20.875000n 0.9  20.975000n 0.9  21.000000n 0.9  21.100000n 0.9  21.125000n 0.9  21.225000n 0.9  21.250000n 0.9  21.350000n 0.9  21.375000n 0.9  21.475000n 0.9  21.500000n 0.9  21.600000n 0.9  21.625000n 0.9  21.725000n 0.9  21.750000n 0.9  21.850000n 0.9  21.875000n 0.9  21.975000n 0.9  22.000000n 0.9  22.100000n 0.9  22.125000n 0.0  22.225000n 0.0  22.250000n 0.0  22.350000n 0.0  22.375000n 0.0  22.475000n 0.0  22.500000n 0.0  22.600000n 0.0  22.625000n 0.0  22.725000n 0.0  22.750000n 0.0  22.850000n 0.0  22.875000n 0.9  22.975000n 0.9  23.000000n 0.9  23.100000n 0.9  23.125000n 0.9  23.225000n 0.9  23.250000n 0.9  23.350000n 0.9  23.375000n 0.9  23.475000n 0.9  23.500000n 0.9  23.600000n 0.9  23.625000n 0.9  23.725000n 0.9  23.750000n 0.9  23.850000n 0.9  23.875000n 0.9  23.975000n 0.9  24.000000n 0.9  24.100000n 0.9  24.125000n 0.9  24.225000n 0.9  24.250000n 0.9  24.350000n 0.9  24.375000n 0.0  24.475000n 0.0  24.500000n 0.0  24.600000n 0.0  24.625000n 0.0  24.725000n 0.0  24.750000n 0.0  24.850000n 0.0  24.875000n 0.0  24.975000n 0.0  25.000000n 0.0  25.100000n 0.0  25.125000n 0.9  25.225000n 0.9  25.250000n 0.9  25.350000n 0.9  25.375000n 0.9  25.475000n 0.9  25.500000n 0.9  25.600000n 0.9  25.625000n 0.9  25.725000n 0.9  25.750000n 0.9  25.850000n 0.9  25.875000n 0.9  25.975000n 0.9  26.000000n 0.9  26.100000n 0.9  26.125000n 0.9  26.225000n 0.9  26.250000n 0.9  26.350000n 0.9  26.375000n 0.9  26.475000n 0.9  26.500000n 0.9  26.600000n 0.9  26.625000n 0.0  26.725000n 0.0  26.750000n 0.0  26.850000n 0.0  26.875000n 0.0  26.975000n 0.0  27.000000n 0.0  27.100000n 0.0  27.125000n 0.0  27.225000n 0.0  27.250000n 0.0  27.350000n 0.0  27.375000n 0.9  27.475000n 0.9  27.500000n 0.9  27.600000n 0.9  27.625000n 0.9  27.725000n 0.9  27.750000n 0.9  27.850000n 0.9  27.875000n 0.9  27.975000n 0.9  28.000000n 0.9  28.100000n 0.9  28.125000n 0.9  28.225000n 0.9  28.250000n 0.9  28.350000n 0.9  28.375000n 0.9  28.475000n 0.9  28.500000n 0.9  28.600000n 0.9  28.625000n 0.9  28.725000n 0.9  28.750000n 0.9  28.850000n 0.9  28.875000n 0.0  28.975000n 0.0  29.000000n 0.0  29.100000n 0.0  29.125000n 0.0  29.225000n 0.0  29.250000n 0.0  29.350000n 0.0  29.375000n 0.0  29.475000n 0.0  29.500000n 0.0  29.600000n 0.0  29.625000n 0.9  29.725000n 0.9  29.750000n 0.9  29.850000n 0.9  29.875000n 0.9  29.975000n 0.9  30.000000n 0.9  30.100000n 0.9  30.125000n 0.9  30.225000n 0.9  30.250000n 0.9 )
V_W20<2> W20<2> W20<1> 0v
V_W20<1> W20<1> 0 PWL(0.000000n 0.0  0.100000n 0.0  0.125000n 0.0  0.225000n 0.0  0.250000n 0.9  0.350000n 0.9  0.375000n 0.9  0.475000n 0.9  0.500000n 0.0  0.600000n 0.0  0.625000n 0.0  0.725000n 0.0  0.750000n 0.0  0.850000n 0.0  0.875000n 0.0  0.975000n 0.0  1.000000n 0.9  1.100000n 0.9  1.125000n 0.9  1.225000n 0.9  1.250000n 0.0  1.350000n 0.0  1.375000n 0.0  1.475000n 0.0  1.500000n 0.0  1.600000n 0.0  1.625000n 0.0  1.725000n 0.0  1.750000n 0.9  1.850000n 0.9  1.875000n 0.9  1.975000n 0.9  2.000000n 0.0  2.100000n 0.0  2.125000n 0.0  2.225000n 0.0  2.250000n 0.0  2.350000n 0.0  2.375000n 0.0  2.475000n 0.0  2.500000n 0.9  2.600000n 0.9  2.625000n 0.9  2.725000n 0.9  2.750000n 0.0  2.850000n 0.0  2.875000n 0.0  2.975000n 0.0  3.000000n 0.0  3.100000n 0.0  3.125000n 0.0  3.225000n 0.0  3.250000n 0.9  3.350000n 0.9  3.375000n 0.9  3.475000n 0.9  3.500000n 0.0  3.600000n 0.0  3.625000n 0.0  3.725000n 0.0  3.750000n 0.0  3.850000n 0.0  3.875000n 0.0  3.975000n 0.0  4.000000n 0.9  4.100000n 0.9  4.125000n 0.9  4.225000n 0.9  4.250000n 0.0  4.350000n 0.0  4.375000n 0.0  4.475000n 0.0  4.500000n 0.0  4.600000n 0.0  4.625000n 0.0  4.725000n 0.0  4.750000n 0.9  4.850000n 0.9  4.875000n 0.9  4.975000n 0.9  5.000000n 0.0  5.100000n 0.0  5.125000n 0.0  5.225000n 0.0  5.250000n 0.0  5.350000n 0.0  5.375000n 0.0  5.475000n 0.0  5.500000n 0.9  5.600000n 0.9  5.625000n 0.9  5.725000n 0.9  5.750000n 0.0  5.850000n 0.0  5.875000n 0.0  5.975000n 0.0  6.000000n 0.0  6.100000n 0.0  6.125000n 0.0  6.225000n 0.0  6.250000n 0.9  6.350000n 0.9  6.375000n 0.9  6.475000n 0.9  6.500000n 0.0  6.600000n 0.0  6.625000n 0.0  6.725000n 0.0  6.750000n 0.0  6.850000n 0.0  6.875000n 0.0  6.975000n 0.0  7.000000n 0.9  7.100000n 0.9  7.125000n 0.9  7.225000n 0.9  7.250000n 0.0  7.350000n 0.0  7.375000n 0.0  7.475000n 0.0  7.500000n 0.0  7.600000n 0.0  7.625000n 0.0  7.725000n 0.0  7.750000n 0.9  7.850000n 0.9  7.875000n 0.9  7.975000n 0.9  8.000000n 0.0  8.100000n 0.0  8.125000n 0.0  8.225000n 0.0  8.250000n 0.0  8.350000n 0.0  8.375000n 0.0  8.475000n 0.0  8.500000n 0.9  8.600000n 0.9  8.625000n 0.9  8.725000n 0.9  8.750000n 0.0  8.850000n 0.0  8.875000n 0.0  8.975000n 0.0  9.000000n 0.0  9.100000n 0.0  9.125000n 0.0  9.225000n 0.0  9.250000n 0.9  9.350000n 0.9  9.375000n 0.9  9.475000n 0.9  9.500000n 0.0  9.600000n 0.0  9.625000n 0.0  9.725000n 0.0  9.750000n 0.0  9.850000n 0.0  9.875000n 0.0  9.975000n 0.0  10.000000n 0.9  10.100000n 0.9  10.125000n 0.9  10.225000n 0.9  10.250000n 0.0  10.350000n 0.0  10.375000n 0.0  10.475000n 0.0  10.500000n 0.0  10.600000n 0.0  10.625000n 0.0  10.725000n 0.0  10.750000n 0.9  10.850000n 0.9  10.875000n 0.9  10.975000n 0.9  11.000000n 0.0  11.100000n 0.0  11.125000n 0.0  11.225000n 0.0  11.250000n 0.0  11.350000n 0.0  11.375000n 0.0  11.475000n 0.0  11.500000n 0.9  11.600000n 0.9  11.625000n 0.9  11.725000n 0.9  11.750000n 0.0  11.850000n 0.0  11.875000n 0.0  11.975000n 0.0  12.000000n 0.0  12.100000n 0.0  12.125000n 0.0  12.225000n 0.0  12.250000n 0.9  12.350000n 0.9  12.375000n 0.9  12.475000n 0.9  12.500000n 0.0  12.600000n 0.0  12.625000n 0.0  12.725000n 0.0  12.750000n 0.0  12.850000n 0.0  12.875000n 0.0  12.975000n 0.0  13.000000n 0.9  13.100000n 0.9  13.125000n 0.9  13.225000n 0.9  13.250000n 0.0  13.350000n 0.0  13.375000n 0.0  13.475000n 0.0  13.500000n 0.0  13.600000n 0.0  13.625000n 0.0  13.725000n 0.0  13.750000n 0.9  13.850000n 0.9  13.875000n 0.9  13.975000n 0.9  14.000000n 0.0  14.100000n 0.0  14.125000n 0.0  14.225000n 0.0  14.250000n 0.0  14.350000n 0.0  14.375000n 0.0  14.475000n 0.0  14.500000n 0.9  14.600000n 0.9  14.625000n 0.9  14.725000n 0.9  14.750000n 0.0  14.850000n 0.0  14.875000n 0.0  14.975000n 0.0  15.000000n 0.0  15.100000n 0.0  15.125000n 0.0  15.225000n 0.0  15.250000n 0.9  15.350000n 0.9  15.375000n 0.9  15.475000n 0.9  15.500000n 0.0  15.600000n 0.0  15.625000n 0.0  15.725000n 0.0  15.750000n 0.0  15.850000n 0.0  15.875000n 0.0  15.975000n 0.0  16.000000n 0.9  16.100000n 0.9  16.125000n 0.9  16.225000n 0.9  16.250000n 0.0  16.350000n 0.0  16.375000n 0.0  16.475000n 0.0  16.500000n 0.0  16.600000n 0.0  16.625000n 0.0  16.725000n 0.0  16.750000n 0.9  16.850000n 0.9  16.875000n 0.9  16.975000n 0.9  17.000000n 0.0  17.100000n 0.0  17.125000n 0.0  17.225000n 0.0  17.250000n 0.0  17.350000n 0.0  17.375000n 0.0  17.475000n 0.0  17.500000n 0.9  17.600000n 0.9  17.625000n 0.9  17.725000n 0.9  17.750000n 0.0  17.850000n 0.0  17.875000n 0.0  17.975000n 0.0  18.000000n 0.0  18.100000n 0.0  18.125000n 0.0  18.225000n 0.0  18.250000n 0.9  18.350000n 0.9  18.375000n 0.9  18.475000n 0.9  18.500000n 0.0  18.600000n 0.0  18.625000n 0.0  18.725000n 0.0  18.750000n 0.0  18.850000n 0.0  18.875000n 0.0  18.975000n 0.0  19.000000n 0.9  19.100000n 0.9  19.125000n 0.9  19.225000n 0.9  19.250000n 0.0  19.350000n 0.0  19.375000n 0.0  19.475000n 0.0  19.500000n 0.0  19.600000n 0.0  19.625000n 0.0  19.725000n 0.0  19.750000n 0.9  19.850000n 0.9  19.875000n 0.9  19.975000n 0.9  20.000000n 0.0  20.100000n 0.0  20.125000n 0.0  20.225000n 0.0  20.250000n 0.0  20.350000n 0.0  20.375000n 0.0  20.475000n 0.0  20.500000n 0.9  20.600000n 0.9  20.625000n 0.9  20.725000n 0.9  20.750000n 0.0  20.850000n 0.0  20.875000n 0.0  20.975000n 0.0  21.000000n 0.0  21.100000n 0.0  21.125000n 0.0  21.225000n 0.0  21.250000n 0.9  21.350000n 0.9  21.375000n 0.9  21.475000n 0.9  21.500000n 0.0  21.600000n 0.0  21.625000n 0.0  21.725000n 0.0  21.750000n 0.0  21.850000n 0.0  21.875000n 0.0  21.975000n 0.0  22.000000n 0.9  22.100000n 0.9  22.125000n 0.9  22.225000n 0.9  22.250000n 0.0  22.350000n 0.0  22.375000n 0.0  22.475000n 0.0  22.500000n 0.0  22.600000n 0.0  22.625000n 0.0  22.725000n 0.0  22.750000n 0.9  22.850000n 0.9  22.875000n 0.9  22.975000n 0.9  23.000000n 0.0  23.100000n 0.0  23.125000n 0.0  23.225000n 0.0  23.250000n 0.0  23.350000n 0.0  23.375000n 0.0  23.475000n 0.0  23.500000n 0.9  23.600000n 0.9  23.625000n 0.9  23.725000n 0.9  23.750000n 0.0  23.850000n 0.0  23.875000n 0.0  23.975000n 0.0  24.000000n 0.0  24.100000n 0.0  24.125000n 0.0  24.225000n 0.0  24.250000n 0.9  24.350000n 0.9  24.375000n 0.9  24.475000n 0.9  24.500000n 0.0  24.600000n 0.0  24.625000n 0.0  24.725000n 0.0  24.750000n 0.0  24.850000n 0.0  24.875000n 0.0  24.975000n 0.0  25.000000n 0.9  25.100000n 0.9  25.125000n 0.9  25.225000n 0.9  25.250000n 0.0  25.350000n 0.0  25.375000n 0.0  25.475000n 0.0  25.500000n 0.0  25.600000n 0.0  25.625000n 0.0  25.725000n 0.0  25.750000n 0.9  25.850000n 0.9  25.875000n 0.9  25.975000n 0.9  26.000000n 0.0  26.100000n 0.0  26.125000n 0.0  26.225000n 0.0  26.250000n 0.0  26.350000n 0.0  26.375000n 0.0  26.475000n 0.0  26.500000n 0.9  26.600000n 0.9  26.625000n 0.9  26.725000n 0.9  26.750000n 0.0  26.850000n 0.0  26.875000n 0.0  26.975000n 0.0  27.000000n 0.0  27.100000n 0.0  27.125000n 0.0  27.225000n 0.0  27.250000n 0.9  27.350000n 0.9  27.375000n 0.9  27.475000n 0.9  27.500000n 0.0  27.600000n 0.0  27.625000n 0.0  27.725000n 0.0  27.750000n 0.0  27.850000n 0.0  27.875000n 0.0  27.975000n 0.0  28.000000n 0.9  28.100000n 0.9  28.125000n 0.9  28.225000n 0.9  28.250000n 0.0  28.350000n 0.0  28.375000n 0.0  28.475000n 0.0  28.500000n 0.0  28.600000n 0.0  28.625000n 0.0  28.725000n 0.0  28.750000n 0.9  28.850000n 0.9  28.875000n 0.9  28.975000n 0.9  29.000000n 0.0  29.100000n 0.0  29.125000n 0.0  29.225000n 0.0  29.250000n 0.0  29.350000n 0.0  29.375000n 0.0  29.475000n 0.0  29.500000n 0.9  29.600000n 0.9  29.625000n 0.9  29.725000n 0.9  29.750000n 0.0  29.850000n 0.0  29.875000n 0.0  29.975000n 0.0  30.000000n 0.0  30.100000n 0.0  30.125000n 0.0  30.225000n 0.0  30.250000n 0.9 )
V_W20<0> W20<0> 0 PWL(0.000000n 0.0  0.100000n 0.0  0.125000n 0.9  0.225000n 0.9  0.250000n 0.9  0.350000n 0.9  0.375000n 0.9  0.475000n 0.9  0.500000n 0.9  0.600000n 0.9  0.625000n 0.0  0.725000n 0.0  0.750000n 0.0  0.850000n 0.0  0.875000n 0.9  0.975000n 0.9  1.000000n 0.9  1.100000n 0.9  1.125000n 0.9  1.225000n 0.9  1.250000n 0.9  1.350000n 0.9  1.375000n 0.0  1.475000n 0.0  1.500000n 0.0  1.600000n 0.0  1.625000n 0.9  1.725000n 0.9  1.750000n 0.9  1.850000n 0.9  1.875000n 0.9  1.975000n 0.9  2.000000n 0.9  2.100000n 0.9  2.125000n 0.0  2.225000n 0.0  2.250000n 0.0  2.350000n 0.0  2.375000n 0.9  2.475000n 0.9  2.500000n 0.9  2.600000n 0.9  2.625000n 0.9  2.725000n 0.9  2.750000n 0.9  2.850000n 0.9  2.875000n 0.0  2.975000n 0.0  3.000000n 0.0  3.100000n 0.0  3.125000n 0.9  3.225000n 0.9  3.250000n 0.9  3.350000n 0.9  3.375000n 0.9  3.475000n 0.9  3.500000n 0.9  3.600000n 0.9  3.625000n 0.0  3.725000n 0.0  3.750000n 0.0  3.850000n 0.0  3.875000n 0.9  3.975000n 0.9  4.000000n 0.9  4.100000n 0.9  4.125000n 0.9  4.225000n 0.9  4.250000n 0.9  4.350000n 0.9  4.375000n 0.0  4.475000n 0.0  4.500000n 0.0  4.600000n 0.0  4.625000n 0.9  4.725000n 0.9  4.750000n 0.9  4.850000n 0.9  4.875000n 0.9  4.975000n 0.9  5.000000n 0.9  5.100000n 0.9  5.125000n 0.0  5.225000n 0.0  5.250000n 0.0  5.350000n 0.0  5.375000n 0.9  5.475000n 0.9  5.500000n 0.9  5.600000n 0.9  5.625000n 0.9  5.725000n 0.9  5.750000n 0.9  5.850000n 0.9  5.875000n 0.0  5.975000n 0.0  6.000000n 0.0  6.100000n 0.0  6.125000n 0.9  6.225000n 0.9  6.250000n 0.9  6.350000n 0.9  6.375000n 0.9  6.475000n 0.9  6.500000n 0.9  6.600000n 0.9  6.625000n 0.0  6.725000n 0.0  6.750000n 0.0  6.850000n 0.0  6.875000n 0.9  6.975000n 0.9  7.000000n 0.9  7.100000n 0.9  7.125000n 0.9  7.225000n 0.9  7.250000n 0.9  7.350000n 0.9  7.375000n 0.0  7.475000n 0.0  7.500000n 0.0  7.600000n 0.0  7.625000n 0.9  7.725000n 0.9  7.750000n 0.9  7.850000n 0.9  7.875000n 0.9  7.975000n 0.9  8.000000n 0.9  8.100000n 0.9  8.125000n 0.0  8.225000n 0.0  8.250000n 0.0  8.350000n 0.0  8.375000n 0.9  8.475000n 0.9  8.500000n 0.9  8.600000n 0.9  8.625000n 0.9  8.725000n 0.9  8.750000n 0.9  8.850000n 0.9  8.875000n 0.0  8.975000n 0.0  9.000000n 0.0  9.100000n 0.0  9.125000n 0.9  9.225000n 0.9  9.250000n 0.9  9.350000n 0.9  9.375000n 0.9  9.475000n 0.9  9.500000n 0.9  9.600000n 0.9  9.625000n 0.0  9.725000n 0.0  9.750000n 0.0  9.850000n 0.0  9.875000n 0.9  9.975000n 0.9  10.000000n 0.9  10.100000n 0.9  10.125000n 0.9  10.225000n 0.9  10.250000n 0.9  10.350000n 0.9  10.375000n 0.0  10.475000n 0.0  10.500000n 0.0  10.600000n 0.0  10.625000n 0.9  10.725000n 0.9  10.750000n 0.9  10.850000n 0.9  10.875000n 0.9  10.975000n 0.9  11.000000n 0.9  11.100000n 0.9  11.125000n 0.0  11.225000n 0.0  11.250000n 0.0  11.350000n 0.0  11.375000n 0.9  11.475000n 0.9  11.500000n 0.9  11.600000n 0.9  11.625000n 0.9  11.725000n 0.9  11.750000n 0.9  11.850000n 0.9  11.875000n 0.0  11.975000n 0.0  12.000000n 0.0  12.100000n 0.0  12.125000n 0.9  12.225000n 0.9  12.250000n 0.9  12.350000n 0.9  12.375000n 0.9  12.475000n 0.9  12.500000n 0.9  12.600000n 0.9  12.625000n 0.0  12.725000n 0.0  12.750000n 0.0  12.850000n 0.0  12.875000n 0.9  12.975000n 0.9  13.000000n 0.9  13.100000n 0.9  13.125000n 0.9  13.225000n 0.9  13.250000n 0.9  13.350000n 0.9  13.375000n 0.0  13.475000n 0.0  13.500000n 0.0  13.600000n 0.0  13.625000n 0.9  13.725000n 0.9  13.750000n 0.9  13.850000n 0.9  13.875000n 0.9  13.975000n 0.9  14.000000n 0.9  14.100000n 0.9  14.125000n 0.0  14.225000n 0.0  14.250000n 0.0  14.350000n 0.0  14.375000n 0.9  14.475000n 0.9  14.500000n 0.9  14.600000n 0.9  14.625000n 0.9  14.725000n 0.9  14.750000n 0.9  14.850000n 0.9  14.875000n 0.0  14.975000n 0.0  15.000000n 0.0  15.100000n 0.0  15.125000n 0.9  15.225000n 0.9  15.250000n 0.9  15.350000n 0.9  15.375000n 0.9  15.475000n 0.9  15.500000n 0.9  15.600000n 0.9  15.625000n 0.0  15.725000n 0.0  15.750000n 0.0  15.850000n 0.0  15.875000n 0.9  15.975000n 0.9  16.000000n 0.9  16.100000n 0.9  16.125000n 0.9  16.225000n 0.9  16.250000n 0.9  16.350000n 0.9  16.375000n 0.0  16.475000n 0.0  16.500000n 0.0  16.600000n 0.0  16.625000n 0.9  16.725000n 0.9  16.750000n 0.9  16.850000n 0.9  16.875000n 0.9  16.975000n 0.9  17.000000n 0.9  17.100000n 0.9  17.125000n 0.0  17.225000n 0.0  17.250000n 0.0  17.350000n 0.0  17.375000n 0.9  17.475000n 0.9  17.500000n 0.9  17.600000n 0.9  17.625000n 0.9  17.725000n 0.9  17.750000n 0.9  17.850000n 0.9  17.875000n 0.0  17.975000n 0.0  18.000000n 0.0  18.100000n 0.0  18.125000n 0.9  18.225000n 0.9  18.250000n 0.9  18.350000n 0.9  18.375000n 0.9  18.475000n 0.9  18.500000n 0.9  18.600000n 0.9  18.625000n 0.0  18.725000n 0.0  18.750000n 0.0  18.850000n 0.0  18.875000n 0.9  18.975000n 0.9  19.000000n 0.9  19.100000n 0.9  19.125000n 0.9  19.225000n 0.9  19.250000n 0.9  19.350000n 0.9  19.375000n 0.0  19.475000n 0.0  19.500000n 0.0  19.600000n 0.0  19.625000n 0.9  19.725000n 0.9  19.750000n 0.9  19.850000n 0.9  19.875000n 0.9  19.975000n 0.9  20.000000n 0.9  20.100000n 0.9  20.125000n 0.0  20.225000n 0.0  20.250000n 0.0  20.350000n 0.0  20.375000n 0.9  20.475000n 0.9  20.500000n 0.9  20.600000n 0.9  20.625000n 0.9  20.725000n 0.9  20.750000n 0.9  20.850000n 0.9  20.875000n 0.0  20.975000n 0.0  21.000000n 0.0  21.100000n 0.0  21.125000n 0.9  21.225000n 0.9  21.250000n 0.9  21.350000n 0.9  21.375000n 0.9  21.475000n 0.9  21.500000n 0.9  21.600000n 0.9  21.625000n 0.0  21.725000n 0.0  21.750000n 0.0  21.850000n 0.0  21.875000n 0.9  21.975000n 0.9  22.000000n 0.9  22.100000n 0.9  22.125000n 0.9  22.225000n 0.9  22.250000n 0.9  22.350000n 0.9  22.375000n 0.0  22.475000n 0.0  22.500000n 0.0  22.600000n 0.0  22.625000n 0.9  22.725000n 0.9  22.750000n 0.9  22.850000n 0.9  22.875000n 0.9  22.975000n 0.9  23.000000n 0.9  23.100000n 0.9  23.125000n 0.0  23.225000n 0.0  23.250000n 0.0  23.350000n 0.0  23.375000n 0.9  23.475000n 0.9  23.500000n 0.9  23.600000n 0.9  23.625000n 0.9  23.725000n 0.9  23.750000n 0.9  23.850000n 0.9  23.875000n 0.0  23.975000n 0.0  24.000000n 0.0  24.100000n 0.0  24.125000n 0.9  24.225000n 0.9  24.250000n 0.9  24.350000n 0.9  24.375000n 0.9  24.475000n 0.9  24.500000n 0.9  24.600000n 0.9  24.625000n 0.0  24.725000n 0.0  24.750000n 0.0  24.850000n 0.0  24.875000n 0.9  24.975000n 0.9  25.000000n 0.9  25.100000n 0.9  25.125000n 0.9  25.225000n 0.9  25.250000n 0.9  25.350000n 0.9  25.375000n 0.0  25.475000n 0.0  25.500000n 0.0  25.600000n 0.0  25.625000n 0.9  25.725000n 0.9  25.750000n 0.9  25.850000n 0.9  25.875000n 0.9  25.975000n 0.9  26.000000n 0.9  26.100000n 0.9  26.125000n 0.0  26.225000n 0.0  26.250000n 0.0  26.350000n 0.0  26.375000n 0.9  26.475000n 0.9  26.500000n 0.9  26.600000n 0.9  26.625000n 0.9  26.725000n 0.9  26.750000n 0.9  26.850000n 0.9  26.875000n 0.0  26.975000n 0.0  27.000000n 0.0  27.100000n 0.0  27.125000n 0.9  27.225000n 0.9  27.250000n 0.9  27.350000n 0.9  27.375000n 0.9  27.475000n 0.9  27.500000n 0.9  27.600000n 0.9  27.625000n 0.0  27.725000n 0.0  27.750000n 0.0  27.850000n 0.0  27.875000n 0.9  27.975000n 0.9  28.000000n 0.9  28.100000n 0.9  28.125000n 0.9  28.225000n 0.9  28.250000n 0.9  28.350000n 0.9  28.375000n 0.0  28.475000n 0.0  28.500000n 0.0  28.600000n 0.0  28.625000n 0.9  28.725000n 0.9  28.750000n 0.9  28.850000n 0.9  28.875000n 0.9  28.975000n 0.9  29.000000n 0.9  29.100000n 0.9  29.125000n 0.0  29.225000n 0.0  29.250000n 0.0  29.350000n 0.0  29.375000n 0.9  29.475000n 0.9  29.500000n 0.9  29.600000n 0.9  29.625000n 0.9  29.725000n 0.9  29.750000n 0.9  29.850000n 0.9  29.875000n 0.0  29.975000n 0.0  30.000000n 0.0  30.100000n 0.0  30.125000n 0.9  30.225000n 0.9  30.250000n 0.9 )
V_Y2 Y2 0 PWL(0.000000n 0.0  0.100000n 0.0  0.125000n 0.0  0.225000n 0.0  0.250000n 0.0  0.350000n 0.0  0.375000n 0.0  0.475000n 0.0  0.500000n 0.0  0.600000n 0.0  0.625000n 0.0  0.725000n 0.0  0.750000n 0.0  0.850000n 0.0  0.875000n 0.0  0.975000n 0.0  1.000000n 0.0  1.100000n 0.0  1.125000n 0.0  1.225000n 0.0  1.250000n 0.0  1.350000n 0.0  1.375000n 0.0  1.475000n 0.0  1.500000n 0.0  1.600000n 0.0  1.625000n 0.0  1.725000n 0.0  1.750000n 0.0  1.850000n 0.0  1.875000n 0.0  1.975000n 0.0  2.000000n 0.0  2.100000n 0.0  2.125000n 0.0  2.225000n 0.0  2.250000n 0.0  2.350000n 0.0  2.375000n 0.0  2.475000n 0.0  2.500000n 0.0  2.600000n 0.0  2.625000n 0.0  2.725000n 0.0  2.750000n 0.0  2.850000n 0.0  2.875000n 0.0  2.975000n 0.0  3.000000n 0.0  3.100000n 0.0  3.125000n 0.0  3.225000n 0.0  3.250000n 0.0  3.350000n 0.0  3.375000n 0.0  3.475000n 0.0  3.500000n 0.0  3.600000n 0.0  3.625000n 0.0  3.725000n 0.0  3.750000n 0.0  3.850000n 0.0  3.875000n 0.0  3.975000n 0.0  4.000000n 0.0  4.100000n 0.0  4.125000n 0.0  4.225000n 0.0  4.250000n 0.0  4.350000n 0.0  4.375000n 0.0  4.475000n 0.0  4.500000n 0.0  4.600000n 0.0  4.625000n 0.0  4.725000n 0.0  4.750000n 0.0  4.850000n 0.0  4.875000n 0.0  4.975000n 0.0  5.000000n 0.0  5.100000n 0.0  5.125000n 0.0  5.225000n 0.0  5.250000n 0.0  5.350000n 0.0  5.375000n 0.0  5.475000n 0.0  5.500000n 0.0  5.600000n 0.0  5.625000n 0.0  5.725000n 0.0  5.750000n 0.0  5.850000n 0.0  5.875000n 0.0  5.975000n 0.0  6.000000n 0.0  6.100000n 0.0  6.125000n 0.0  6.225000n 0.0  6.250000n 0.0  6.350000n 0.0  6.375000n 0.0  6.475000n 0.0  6.500000n 0.0  6.600000n 0.0  6.625000n 0.0  6.725000n 0.0  6.750000n 0.0  6.850000n 0.0  6.875000n 0.0  6.975000n 0.0  7.000000n 0.0  7.100000n 0.0  7.125000n 0.0  7.225000n 0.0  7.250000n 0.0  7.350000n 0.0  7.375000n 0.0  7.475000n 0.0  7.500000n 0.0  7.600000n 0.0  7.625000n 0.0  7.725000n 0.0  7.750000n 0.0  7.850000n 0.0  7.875000n 0.0  7.975000n 0.0  8.000000n 0.0  8.100000n 0.0  8.125000n 0.0  8.225000n 0.0  8.250000n 0.0  8.350000n 0.0  8.375000n 0.0  8.475000n 0.0  8.500000n 0.0  8.600000n 0.0  8.625000n 0.0  8.725000n 0.0  8.750000n 0.0  8.850000n 0.0  8.875000n 0.0  8.975000n 0.0  9.000000n 0.0  9.100000n 0.0  9.125000n 0.0  9.225000n 0.0  9.250000n 0.0  9.350000n 0.0  9.375000n 0.0  9.475000n 0.0  9.500000n 0.0  9.600000n 0.0  9.625000n 0.0  9.725000n 0.0  9.750000n 0.0  9.850000n 0.0  9.875000n 0.0  9.975000n 0.0  10.000000n 0.0  10.100000n 0.0  10.125000n 0.0  10.225000n 0.0  10.250000n 0.0  10.350000n 0.0  10.375000n 0.0  10.475000n 0.0  10.500000n 0.0  10.600000n 0.0  10.625000n 0.0  10.725000n 0.0  10.750000n 0.0  10.850000n 0.0  10.875000n 0.0  10.975000n 0.0  11.000000n 0.0  11.100000n 0.0  11.125000n 0.0  11.225000n 0.0  11.250000n 0.0  11.350000n 0.0  11.375000n 0.0  11.475000n 0.0  11.500000n 0.0  11.600000n 0.0  11.625000n 0.0  11.725000n 0.0  11.750000n 0.0  11.850000n 0.0  11.875000n 0.0  11.975000n 0.0  12.000000n 0.0  12.100000n 0.0  12.125000n 0.0  12.225000n 0.0  12.250000n 0.0  12.350000n 0.0  12.375000n 0.0  12.475000n 0.0  12.500000n 0.0  12.600000n 0.0  12.625000n 0.0  12.725000n 0.0  12.750000n 0.0  12.850000n 0.0  12.875000n 0.0  12.975000n 0.0  13.000000n 0.0  13.100000n 0.0  13.125000n 0.0  13.225000n 0.0  13.250000n 0.0  13.350000n 0.0  13.375000n 0.0  13.475000n 0.0  13.500000n 0.0  13.600000n 0.0  13.625000n 0.0  13.725000n 0.0  13.750000n 0.0  13.850000n 0.0  13.875000n 0.0  13.975000n 0.0  14.000000n 0.0  14.100000n 0.0  14.125000n 0.0  14.225000n 0.0  14.250000n 0.0  14.350000n 0.0  14.375000n 0.0  14.475000n 0.0  14.500000n 0.0  14.600000n 0.0  14.625000n 0.0  14.725000n 0.0  14.750000n 0.0  14.850000n 0.0  14.875000n 0.0  14.975000n 0.0  15.000000n 0.0  15.100000n 0.0  15.125000n 0.0  15.225000n 0.0  15.250000n 0.0  15.350000n 0.0  15.375000n 0.0  15.475000n 0.0  15.500000n 0.0  15.600000n 0.0  15.625000n 0.0  15.725000n 0.0  15.750000n 0.0  15.850000n 0.0  15.875000n 0.0  15.975000n 0.0  16.000000n 0.0  16.100000n 0.0  16.125000n 0.0  16.225000n 0.0  16.250000n 0.0  16.350000n 0.0  16.375000n 0.0  16.475000n 0.0  16.500000n 0.0  16.600000n 0.0  16.625000n 0.0  16.725000n 0.0  16.750000n 0.0  16.850000n 0.0  16.875000n 0.0  16.975000n 0.0  17.000000n 0.0  17.100000n 0.0  17.125000n 0.0  17.225000n 0.0  17.250000n 0.0  17.350000n 0.0  17.375000n 0.0  17.475000n 0.0  17.500000n 0.0  17.600000n 0.0  17.625000n 0.0  17.725000n 0.0  17.750000n 0.0  17.850000n 0.0  17.875000n 0.0  17.975000n 0.0  18.000000n 0.0  18.100000n 0.0  18.125000n 0.0  18.225000n 0.0  18.250000n 0.0  18.350000n 0.0  18.375000n 0.0  18.475000n 0.0  18.500000n 0.0  18.600000n 0.0  18.625000n 0.0  18.725000n 0.0  18.750000n 0.0  18.850000n 0.0  18.875000n 0.0  18.975000n 0.0  19.000000n 0.0  19.100000n 0.0  19.125000n 0.0  19.225000n 0.0  19.250000n 0.0  19.350000n 0.0  19.375000n 0.0  19.475000n 0.0  19.500000n 0.0  19.600000n 0.0  19.625000n 0.0  19.725000n 0.0  19.750000n 0.0  19.850000n 0.0  19.875000n 0.0  19.975000n 0.0  20.000000n 0.0  20.100000n 0.0  20.125000n 0.0  20.225000n 0.0  20.250000n 0.0  20.350000n 0.0  20.375000n 0.0  20.475000n 0.0  20.500000n 0.0  20.600000n 0.0  20.625000n 0.0  20.725000n 0.0  20.750000n 0.0  20.850000n 0.0  20.875000n 0.0  20.975000n 0.0  21.000000n 0.0  21.100000n 0.0  21.125000n 0.0  21.225000n 0.0  21.250000n 0.0  21.350000n 0.0  21.375000n 0.0  21.475000n 0.0  21.500000n 0.0  21.600000n 0.0  21.625000n 0.0  21.725000n 0.0  21.750000n 0.0  21.850000n 0.0  21.875000n 0.0  21.975000n 0.0  22.000000n 0.0  22.100000n 0.0  22.125000n 0.0  22.225000n 0.0  22.250000n 0.0  22.350000n 0.0  22.375000n 0.0  22.475000n 0.0  22.500000n 0.0  22.600000n 0.0  22.625000n 0.0  22.725000n 0.0  22.750000n 0.0  22.850000n 0.0  22.875000n 0.0  22.975000n 0.0  23.000000n 0.0  23.100000n 0.0  23.125000n 0.0  23.225000n 0.0  23.250000n 0.0  23.350000n 0.0  23.375000n 0.0  23.475000n 0.0  23.500000n 0.0  23.600000n 0.0  23.625000n 0.0  23.725000n 0.0  23.750000n 0.0  23.850000n 0.0  23.875000n 0.0  23.975000n 0.0  24.000000n 0.0  24.100000n 0.0  24.125000n 0.0  24.225000n 0.0  24.250000n 0.0  24.350000n 0.0  24.375000n 0.0  24.475000n 0.0  24.500000n 0.0  24.600000n 0.0  24.625000n 0.0  24.725000n 0.0  24.750000n 0.0  24.850000n 0.0  24.875000n 0.0  24.975000n 0.0  25.000000n 0.0  25.100000n 0.0  25.125000n 0.0  25.225000n 0.0  25.250000n 0.0  25.350000n 0.0  25.375000n 0.0  25.475000n 0.0  25.500000n 0.0  25.600000n 0.0  25.625000n 0.0  25.725000n 0.0  25.750000n 0.0  25.850000n 0.0  25.875000n 0.0  25.975000n 0.0  26.000000n 0.0  26.100000n 0.0  26.125000n 0.0  26.225000n 0.0  26.250000n 0.0  26.350000n 0.0  26.375000n 0.0  26.475000n 0.0  26.500000n 0.0  26.600000n 0.0  26.625000n 0.0  26.725000n 0.0  26.750000n 0.0  26.850000n 0.0  26.875000n 0.0  26.975000n 0.0  27.000000n 0.0  27.100000n 0.0  27.125000n 0.0  27.225000n 0.0  27.250000n 0.0  27.350000n 0.0  27.375000n 0.0  27.475000n 0.0  27.500000n 0.0  27.600000n 0.0  27.625000n 0.0  27.725000n 0.0  27.750000n 0.0  27.850000n 0.0  27.875000n 0.0  27.975000n 0.0  28.000000n 0.0  28.100000n 0.0  28.125000n 0.0  28.225000n 0.0  28.250000n 0.0  28.350000n 0.0  28.375000n 0.0  28.475000n 0.0  28.500000n 0.0  28.600000n 0.0  28.625000n 0.0  28.725000n 0.0  28.750000n 0.0  28.850000n 0.0  28.875000n 0.0  28.975000n 0.0  29.000000n 0.0  29.100000n 0.0  29.125000n 0.0  29.225000n 0.0  29.250000n 0.0  29.350000n 0.0  29.375000n 0.0  29.475000n 0.0  29.500000n 0.0  29.600000n 0.0  29.625000n 0.0  29.725000n 0.0  29.750000n 0.0  29.850000n 0.0  29.875000n 0.0  29.975000n 0.0  30.000000n 0.0  30.100000n 0.0  30.125000n 0.0  30.225000n 0.0  30.250000n 0.0 )
V_Y1 Y1 0 PWL(0.000000n 0.0  0.100000n 0.0  0.125000n 0.0  0.225000n 0.0  0.250000n 0.0  0.350000n 0.0  0.375000n 0.0  0.475000n 0.0  0.500000n 0.0  0.600000n 0.0  0.625000n 0.0  0.725000n 0.0  0.750000n 0.0  0.850000n 0.0  0.875000n 0.0  0.975000n 0.0  1.000000n 0.0  1.100000n 0.0  1.125000n 0.0  1.225000n 0.0  1.250000n 0.0  1.350000n 0.0  1.375000n 0.0  1.475000n 0.0  1.500000n 0.0  1.600000n 0.0  1.625000n 0.0  1.725000n 0.0  1.750000n 0.0  1.850000n 0.0  1.875000n 0.0  1.975000n 0.0  2.000000n 0.0  2.100000n 0.0  2.125000n 0.0  2.225000n 0.0  2.250000n 0.0  2.350000n 0.0  2.375000n 0.0  2.475000n 0.0  2.500000n 0.0  2.600000n 0.0  2.625000n 0.0  2.725000n 0.0  2.750000n 0.0  2.850000n 0.0  2.875000n 0.0  2.975000n 0.0  3.000000n 0.0  3.100000n 0.0  3.125000n 0.0  3.225000n 0.0  3.250000n 0.0  3.350000n 0.0  3.375000n 0.0  3.475000n 0.0  3.500000n 0.0  3.600000n 0.0  3.625000n 0.0  3.725000n 0.0  3.750000n 0.0  3.850000n 0.0  3.875000n 0.9  3.975000n 0.9  4.000000n 0.0  4.100000n 0.0  4.125000n 0.0  4.225000n 0.0  4.250000n 0.0  4.350000n 0.0  4.375000n 0.0  4.475000n 0.0  4.500000n 0.0  4.600000n 0.0  4.625000n 0.0  4.725000n 0.0  4.750000n 0.0  4.850000n 0.0  4.875000n 0.0  4.975000n 0.0  5.000000n 0.9  5.100000n 0.9  5.125000n 0.0  5.225000n 0.0  5.250000n 0.0  5.350000n 0.0  5.375000n 0.0  5.475000n 0.0  5.500000n 0.0  5.600000n 0.0  5.625000n 0.0  5.725000n 0.0  5.750000n 0.0  5.850000n 0.0  5.875000n 0.0  5.975000n 0.0  6.000000n 0.0  6.100000n 0.0  6.125000n 0.9  6.225000n 0.9  6.250000n 0.0  6.350000n 0.0  6.375000n 0.0  6.475000n 0.0  6.500000n 0.0  6.600000n 0.0  6.625000n 0.0  6.725000n 0.0  6.750000n 0.0  6.850000n 0.0  6.875000n 0.0  6.975000n 0.0  7.000000n 0.0  7.100000n 0.0  7.125000n 0.0  7.225000n 0.0  7.250000n 0.0  7.350000n 0.0  7.375000n 0.0  7.475000n 0.0  7.500000n 0.0  7.600000n 0.0  7.625000n 0.9  7.725000n 0.9  7.750000n 0.0  7.850000n 0.0  7.875000n 0.0  7.975000n 0.0  8.000000n 0.9  8.100000n 0.9  8.125000n 0.0  8.225000n 0.0  8.250000n 0.0  8.350000n 0.0  8.375000n 0.0  8.475000n 0.0  8.500000n 0.0  8.600000n 0.0  8.625000n 0.0  8.725000n 0.0  8.750000n 0.0  8.850000n 0.0  8.875000n 0.0  8.975000n 0.0  9.000000n 0.0  9.100000n 0.0  9.125000n 0.0  9.225000n 0.0  9.250000n 0.0  9.350000n 0.0  9.375000n 0.0  9.475000n 0.0  9.500000n 0.0  9.600000n 0.0  9.625000n 0.0  9.725000n 0.0  9.750000n 0.0  9.850000n 0.0  9.875000n 0.9  9.975000n 0.9  10.000000n 0.0  10.100000n 0.0  10.125000n 0.0  10.225000n 0.0  10.250000n 0.0  10.350000n 0.0  10.375000n 0.0  10.475000n 0.0  10.500000n 0.0  10.600000n 0.0  10.625000n 0.0  10.725000n 0.0  10.750000n 0.0  10.850000n 0.0  10.875000n 0.0  10.975000n 0.0  11.000000n 0.0  11.100000n 0.0  11.125000n 0.0  11.225000n 0.0  11.250000n 0.0  11.350000n 0.0  11.375000n 0.9  11.475000n 0.9  11.500000n 0.0  11.600000n 0.0  11.625000n 0.0  11.725000n 0.0  11.750000n 0.0  11.850000n 0.0  11.875000n 0.0  11.975000n 0.0  12.000000n 0.9  12.100000n 0.9  12.125000n 0.9  12.225000n 0.9  12.250000n 0.0  12.350000n 0.0  12.375000n 0.0  12.475000n 0.0  12.500000n 0.9  12.600000n 0.9  12.625000n 0.0  12.725000n 0.0  12.750000n 0.0  12.850000n 0.0  12.875000n 0.0  12.975000n 0.0  13.000000n 0.0  13.100000n 0.0  13.125000n 0.0  13.225000n 0.0  13.250000n 0.0  13.350000n 0.0  13.375000n 0.0  13.475000n 0.0  13.500000n 0.0  13.600000n 0.0  13.625000n 0.0  13.725000n 0.0  13.750000n 0.0  13.850000n 0.0  13.875000n 0.0  13.975000n 0.0  14.000000n 0.9  14.100000n 0.9  14.125000n 0.0  14.225000n 0.0  14.250000n 0.0  14.350000n 0.0  14.375000n 0.0  14.475000n 0.0  14.500000n 0.0  14.600000n 0.0  14.625000n 0.0  14.725000n 0.0  14.750000n 0.0  14.850000n 0.0  14.875000n 0.0  14.975000n 0.0  15.000000n 0.9  15.100000n 0.9  15.125000n 0.9  15.225000n 0.9  15.250000n 0.0  15.350000n 0.0  15.375000n 0.0  15.475000n 0.0  15.500000n 0.9  15.600000n 0.9  15.625000n 0.0  15.725000n 0.0  15.750000n 0.0  15.850000n 0.0  15.875000n 0.0  15.975000n 0.0  16.000000n 0.0  16.100000n 0.0  16.125000n 0.0  16.225000n 0.0  16.250000n 0.0  16.350000n 0.0  16.375000n 0.0  16.475000n 0.0  16.500000n 0.0  16.600000n 0.0  16.625000n 0.0  16.725000n 0.0  16.750000n 0.0  16.850000n 0.0  16.875000n 0.0  16.975000n 0.0  17.000000n 0.0  17.100000n 0.0  17.125000n 0.0  17.225000n 0.0  17.250000n 0.0  17.350000n 0.0  17.375000n 0.0  17.475000n 0.0  17.500000n 0.0  17.600000n 0.0  17.625000n 0.0  17.725000n 0.0  17.750000n 0.0  17.850000n 0.0  17.875000n 0.0  17.975000n 0.0  18.000000n 0.0  18.100000n 0.0  18.125000n 0.9  18.225000n 0.9  18.250000n 0.0  18.350000n 0.0  18.375000n 0.0  18.475000n 0.0  18.500000n 0.9  18.600000n 0.9  18.625000n 0.0  18.725000n 0.0  18.750000n 0.0  18.850000n 0.0  18.875000n 0.9  18.975000n 0.9  19.000000n 0.0  19.100000n 0.0  19.125000n 0.0  19.225000n 0.0  19.250000n 0.0  19.350000n 0.0  19.375000n 0.0  19.475000n 0.0  19.500000n 0.0  19.600000n 0.0  19.625000n 0.0  19.725000n 0.0  19.750000n 0.0  19.850000n 0.0  19.875000n 0.0  19.975000n 0.0  20.000000n 0.0  20.100000n 0.0  20.125000n 0.0  20.225000n 0.0  20.250000n 0.0  20.350000n 0.0  20.375000n 0.0  20.475000n 0.0  20.500000n 0.0  20.600000n 0.0  20.625000n 0.0  20.725000n 0.0  20.750000n 0.0  20.850000n 0.0  20.875000n 0.0  20.975000n 0.0  21.000000n 0.0  21.100000n 0.0  21.125000n 0.0  21.225000n 0.0  21.250000n 0.0  21.350000n 0.0  21.375000n 0.0  21.475000n 0.0  21.500000n 0.0  21.600000n 0.0  21.625000n 0.0  21.725000n 0.0  21.750000n 0.0  21.850000n 0.0  21.875000n 0.0  21.975000n 0.0  22.000000n 0.0  22.100000n 0.0  22.125000n 0.0  22.225000n 0.0  22.250000n 0.0  22.350000n 0.0  22.375000n 0.0  22.475000n 0.0  22.500000n 0.0  22.600000n 0.0  22.625000n 0.9  22.725000n 0.9  22.750000n 0.0  22.850000n 0.0  22.875000n 0.0  22.975000n 0.0  23.000000n 0.9  23.100000n 0.9  23.125000n 0.0  23.225000n 0.0  23.250000n 0.0  23.350000n 0.0  23.375000n 0.9  23.475000n 0.9  23.500000n 0.0  23.600000n 0.0  23.625000n 0.0  23.725000n 0.0  23.750000n 0.0  23.850000n 0.0  23.875000n 0.0  23.975000n 0.0  24.000000n 0.9  24.100000n 0.9  24.125000n 0.9  24.225000n 0.9  24.250000n 0.0  24.350000n 0.0  24.375000n 0.0  24.475000n 0.0  24.500000n 0.9  24.600000n 0.9  24.625000n 0.0  24.725000n 0.0  24.750000n 0.0  24.850000n 0.0  24.875000n 0.0  24.975000n 0.0  25.000000n 0.0  25.100000n 0.0  25.125000n 0.0  25.225000n 0.0  25.250000n 0.0  25.350000n 0.0  25.375000n 0.0  25.475000n 0.0  25.500000n 0.0  25.600000n 0.0  25.625000n 0.0  25.725000n 0.0  25.750000n 0.0  25.850000n 0.0  25.875000n 0.0  25.975000n 0.0  26.000000n 0.0  26.100000n 0.0  26.125000n 0.0  26.225000n 0.0  26.250000n 0.0  26.350000n 0.0  26.375000n 0.9  26.475000n 0.9  26.500000n 0.0  26.600000n 0.0  26.625000n 0.0  26.725000n 0.0  26.750000n 0.0  26.850000n 0.0  26.875000n 0.0  26.975000n 0.0  27.000000n 0.0  27.100000n 0.0  27.125000n 0.0  27.225000n 0.0  27.250000n 0.0  27.350000n 0.0  27.375000n 0.0  27.475000n 0.0  27.500000n 0.0  27.600000n 0.0  27.625000n 0.0  27.725000n 0.0  27.750000n 0.0  27.850000n 0.0  27.875000n 0.9  27.975000n 0.9  28.000000n 0.0  28.100000n 0.0  28.125000n 0.0  28.225000n 0.0  28.250000n 0.0  28.350000n 0.0  28.375000n 0.0  28.475000n 0.0  28.500000n 0.0  28.600000n 0.0  28.625000n 0.0  28.725000n 0.0  28.750000n 0.0  28.850000n 0.0  28.875000n 0.0  28.975000n 0.0  29.000000n 0.0  29.100000n 0.0  29.125000n 0.0  29.225000n 0.0  29.250000n 0.0  29.350000n 0.0  29.375000n 0.9  29.475000n 0.9  29.500000n 0.0  29.600000n 0.0  29.625000n 0.0  29.725000n 0.0  29.750000n 0.0  29.850000n 0.0  29.875000n 0.0  29.975000n 0.0  30.000000n 0.9  30.100000n 0.9  30.125000n 0.9  30.225000n 0.9  30.250000n 0.0 )
V_Y0 Y0 0 PWL(0.000000n 0.0  0.100000n 0.0  0.125000n 0.9  0.225000n 0.9  0.250000n 0.0  0.350000n 0.0  0.375000n 0.0  0.475000n 0.0  0.500000n 0.9  0.600000n 0.9  0.625000n 0.0  0.725000n 0.0  0.750000n 0.0  0.850000n 0.0  0.875000n 0.9  0.975000n 0.9  1.000000n 0.0  1.100000n 0.0  1.125000n 0.0  1.225000n 0.0  1.250000n 0.9  1.350000n 0.9  1.375000n 0.0  1.475000n 0.0  1.500000n 0.0  1.600000n 0.0  1.625000n 0.9  1.725000n 0.9  1.750000n 0.0  1.850000n 0.0  1.875000n 0.0  1.975000n 0.0  2.000000n 0.9  2.100000n 0.9  2.125000n 0.0  2.225000n 0.0  2.250000n 0.0  2.350000n 0.0  2.375000n 0.9  2.475000n 0.9  2.500000n 0.0  2.600000n 0.0  2.625000n 0.0  2.725000n 0.0  2.750000n 0.9  2.850000n 0.9  2.875000n 0.0  2.975000n 0.0  3.000000n 0.0  3.100000n 0.0  3.125000n 0.9  3.225000n 0.9  3.250000n 0.0  3.350000n 0.0  3.375000n 0.0  3.475000n 0.0  3.500000n 0.0  3.600000n 0.0  3.625000n 0.0  3.725000n 0.0  3.750000n 0.9  3.850000n 0.9  3.875000n 0.0  3.975000n 0.0  4.000000n 0.0  4.100000n 0.0  4.125000n 0.0  4.225000n 0.0  4.250000n 0.9  4.350000n 0.9  4.375000n 0.0  4.475000n 0.0  4.500000n 0.0  4.600000n 0.0  4.625000n 0.9  4.725000n 0.9  4.750000n 0.0  4.850000n 0.0  4.875000n 0.0  4.975000n 0.0  5.000000n 0.0  5.100000n 0.0  5.125000n 0.9  5.225000n 0.9  5.250000n 0.0  5.350000n 0.0  5.375000n 0.0  5.475000n 0.0  5.500000n 0.0  5.600000n 0.0  5.625000n 0.0  5.725000n 0.0  5.750000n 0.0  5.850000n 0.0  5.875000n 0.0  5.975000n 0.0  6.000000n 0.9  6.100000n 0.9  6.125000n 0.0  6.225000n 0.0  6.250000n 0.0  6.350000n 0.0  6.375000n 0.0  6.475000n 0.0  6.500000n 0.9  6.600000n 0.9  6.625000n 0.0  6.725000n 0.0  6.750000n 0.0  6.850000n 0.0  6.875000n 0.9  6.975000n 0.9  7.000000n 0.0  7.100000n 0.0  7.125000n 0.0  7.225000n 0.0  7.250000n 0.0  7.350000n 0.0  7.375000n 0.0  7.475000n 0.0  7.500000n 0.9  7.600000n 0.9  7.625000n 0.0  7.725000n 0.0  7.750000n 0.0  7.850000n 0.0  7.875000n 0.0  7.975000n 0.0  8.000000n 0.0  8.100000n 0.0  8.125000n 0.9  8.225000n 0.9  8.250000n 0.0  8.350000n 0.0  8.375000n 0.0  8.475000n 0.0  8.500000n 0.0  8.600000n 0.0  8.625000n 0.0  8.725000n 0.0  8.750000n 0.9  8.850000n 0.9  8.875000n 0.0  8.975000n 0.0  9.000000n 0.0  9.100000n 0.0  9.125000n 0.9  9.225000n 0.9  9.250000n 0.0  9.350000n 0.0  9.375000n 0.0  9.475000n 0.0  9.500000n 0.0  9.600000n 0.0  9.625000n 0.0  9.725000n 0.0  9.750000n 0.9  9.850000n 0.9  9.875000n 0.0  9.975000n 0.0  10.000000n 0.0  10.100000n 0.0  10.125000n 0.0  10.225000n 0.0  10.250000n 0.9  10.350000n 0.9  10.375000n 0.0  10.475000n 0.0  10.500000n 0.0  10.600000n 0.0  10.625000n 0.0  10.725000n 0.0  10.750000n 0.0  10.850000n 0.0  10.875000n 0.0  10.975000n 0.0  11.000000n 0.0  11.100000n 0.0  11.125000n 0.0  11.225000n 0.0  11.250000n 0.9  11.350000n 0.9  11.375000n 0.0  11.475000n 0.0  11.500000n 0.0  11.600000n 0.0  11.625000n 0.0  11.725000n 0.0  11.750000n 0.9  11.850000n 0.9  11.875000n 0.0  11.975000n 0.0  12.000000n 0.0  12.100000n 0.0  12.125000n 0.9  12.225000n 0.9  12.250000n 0.9  12.350000n 0.9  12.375000n 0.0  12.475000n 0.0  12.500000n 0.0  12.600000n 0.0  12.625000n 0.9  12.725000n 0.9  12.750000n 0.0  12.850000n 0.0  12.875000n 0.0  12.975000n 0.0  13.000000n 0.0  13.100000n 0.0  13.125000n 0.0  13.225000n 0.0  13.250000n 0.9  13.350000n 0.9  13.375000n 0.0  13.475000n 0.0  13.500000n 0.0  13.600000n 0.0  13.625000n 0.9  13.725000n 0.9  13.750000n 0.0  13.850000n 0.0  13.875000n 0.0  13.975000n 0.0  14.000000n 0.0  14.100000n 0.0  14.125000n 0.9  14.225000n 0.9  14.250000n 0.0  14.350000n 0.0  14.375000n 0.0  14.475000n 0.0  14.500000n 0.0  14.600000n 0.0  14.625000n 0.0  14.725000n 0.0  14.750000n 0.9  14.850000n 0.9  14.875000n 0.0  14.975000n 0.0  15.000000n 0.0  15.100000n 0.0  15.125000n 0.9  15.225000n 0.9  15.250000n 0.9  15.350000n 0.9  15.375000n 0.0  15.475000n 0.0  15.500000n 0.0  15.600000n 0.0  15.625000n 0.9  15.725000n 0.9  15.750000n 0.0  15.850000n 0.0  15.875000n 0.0  15.975000n 0.0  16.000000n 0.0  16.100000n 0.0  16.125000n 0.0  16.225000n 0.0  16.250000n 0.9  16.350000n 0.9  16.375000n 0.0  16.475000n 0.0  16.500000n 0.0  16.600000n 0.0  16.625000n 0.0  16.725000n 0.0  16.750000n 0.0  16.850000n 0.0  16.875000n 0.0  16.975000n 0.0  17.000000n 0.0  17.100000n 0.0  17.125000n 0.0  17.225000n 0.0  17.250000n 0.0  17.350000n 0.0  17.375000n 0.0  17.475000n 0.0  17.500000n 0.0  17.600000n 0.0  17.625000n 0.0  17.725000n 0.0  17.750000n 0.0  17.850000n 0.0  17.875000n 0.0  17.975000n 0.0  18.000000n 0.9  18.100000n 0.9  18.125000n 0.0  18.225000n 0.0  18.250000n 0.0  18.350000n 0.0  18.375000n 0.0  18.475000n 0.0  18.500000n 0.0  18.600000n 0.0  18.625000n 0.9  18.725000n 0.9  18.750000n 0.9  18.850000n 0.9  18.875000n 0.0  18.975000n 0.0  19.000000n 0.0  19.100000n 0.0  19.125000n 0.0  19.225000n 0.0  19.250000n 0.9  19.350000n 0.9  19.375000n 0.0  19.475000n 0.0  19.500000n 0.0  19.600000n 0.0  19.625000n 0.9  19.725000n 0.9  19.750000n 0.0  19.850000n 0.0  19.875000n 0.0  19.975000n 0.0  20.000000n 0.9  20.100000n 0.9  20.125000n 0.0  20.225000n 0.0  20.250000n 0.0  20.350000n 0.0  20.375000n 0.9  20.475000n 0.9  20.500000n 0.0  20.600000n 0.0  20.625000n 0.0  20.725000n 0.0  20.750000n 0.9  20.850000n 0.9  20.875000n 0.0  20.975000n 0.0  21.000000n 0.0  21.100000n 0.0  21.125000n 0.9  21.225000n 0.9  21.250000n 0.0  21.350000n 0.0  21.375000n 0.0  21.475000n 0.0  21.500000n 0.0  21.600000n 0.0  21.625000n 0.0  21.725000n 0.0  21.750000n 0.0  21.850000n 0.0  21.875000n 0.0  21.975000n 0.0  22.000000n 0.0  22.100000n 0.0  22.125000n 0.0  22.225000n 0.0  22.250000n 0.0  22.350000n 0.0  22.375000n 0.0  22.475000n 0.0  22.500000n 0.9  22.600000n 0.9  22.625000n 0.0  22.725000n 0.0  22.750000n 0.0  22.850000n 0.0  22.875000n 0.0  22.975000n 0.0  23.000000n 0.0  23.100000n 0.0  23.125000n 0.9  23.225000n 0.9  23.250000n 0.9  23.350000n 0.9  23.375000n 0.0  23.475000n 0.0  23.500000n 0.0  23.600000n 0.0  23.625000n 0.0  23.725000n 0.0  23.750000n 0.9  23.850000n 0.9  23.875000n 0.0  23.975000n 0.0  24.000000n 0.0  24.100000n 0.0  24.125000n 0.9  24.225000n 0.9  24.250000n 0.9  24.350000n 0.9  24.375000n 0.0  24.475000n 0.0  24.500000n 0.0  24.600000n 0.0  24.625000n 0.9  24.725000n 0.9  24.750000n 0.0  24.850000n 0.0  24.875000n 0.0  24.975000n 0.0  25.000000n 0.0  25.100000n 0.0  25.125000n 0.0  25.225000n 0.0  25.250000n 0.9  25.350000n 0.9  25.375000n 0.0  25.475000n 0.0  25.500000n 0.0  25.600000n 0.0  25.625000n 0.0  25.725000n 0.0  25.750000n 0.0  25.850000n 0.0  25.875000n 0.0  25.975000n 0.0  26.000000n 0.0  26.100000n 0.0  26.125000n 0.0  26.225000n 0.0  26.250000n 0.9  26.350000n 0.9  26.375000n 0.0  26.475000n 0.0  26.500000n 0.0  26.600000n 0.0  26.625000n 0.0  26.725000n 0.0  26.750000n 0.9  26.850000n 0.9  26.875000n 0.0  26.975000n 0.0  27.000000n 0.0  27.100000n 0.0  27.125000n 0.9  27.225000n 0.9  27.250000n 0.0  27.350000n 0.0  27.375000n 0.0  27.475000n 0.0  27.500000n 0.0  27.600000n 0.0  27.625000n 0.0  27.725000n 0.0  27.750000n 0.9  27.850000n 0.9  27.875000n 0.0  27.975000n 0.0  28.000000n 0.0  28.100000n 0.0  28.125000n 0.0  28.225000n 0.0  28.250000n 0.9  28.350000n 0.9  28.375000n 0.0  28.475000n 0.0  28.500000n 0.0  28.600000n 0.0  28.625000n 0.0  28.725000n 0.0  28.750000n 0.0  28.850000n 0.0  28.875000n 0.0  28.975000n 0.0  29.000000n 0.0  29.100000n 0.0  29.125000n 0.0  29.225000n 0.0  29.250000n 0.9  29.350000n 0.9  29.375000n 0.0  29.475000n 0.0  29.500000n 0.0  29.600000n 0.0  29.625000n 0.0  29.725000n 0.0  29.750000n 0.9  29.850000n 0.9  29.875000n 0.0  29.975000n 0.0  30.000000n 0.0  30.100000n 0.0  30.125000n 0.9  30.225000n 0.9  30.250000n 0.9 )


* Set fanout manually or by instantiating four other inverters
* cout out vss! 100f

* Transient analysis
.TRAN 5p 30.5n

